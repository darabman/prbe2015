-- =============================================================================================================
-- *
-- * Copyright (c) University of York
-- *
-- * File Name: internal_rom_64K.vhd
-- *
-- * Version: V1.0
-- *
-- * Release Date:
-- *
-- * Author(s): M.Freeman
-- *
-- * Description: Read Only Memory based on blockRams 
-- *
-- * Change History:  $Author: $
-- *                  $Date: $
-- *                  $Revision: $
-- *
-- * Conditions of Use: THIS CODE IS COPYRIGHT AND IS SUPPLIED "AS IS" WITHOUT WARRANTY OF ANY KIND, INCLUDING,
-- *                    BUT NOT LIMITED TO, ANY IMPLIED WARRANTY OF MERCHANTABILITY AND FITNESS FOR A
-- *                    PARTICULAR PURPOSE.
-- *
-- * Notes:
-- *
-- =============================================================================================================

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

LIBRARY UNISIM;
USE UNISIM.vcomponents.ALL;

LIBRARY work;
USE work.internal_rom_64K_pkg.ALL ;

ENTITY internal_rom_64K IS 
PORT (
  clk_i : IN STD_LOGIC;
  rst_i : IN STD_LOGIC;
  adr_i : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
  dat_o : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
  stb_i : IN STD_LOGIC; 
  cyc_i : IN STD_LOGIC; 
  ack_o : OUT STD_LOGIC );  
END internal_rom_64K;

ARCHITECTURE internal_rom_64K_arch OF internal_rom_64K IS 

  --
  -- components
  --

  COMPONENT RAMB16_S9
  GENERIC(
    INIT_00 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
    INIT_01 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
    INIT_02 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
    INIT_03 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
    INIT_04 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
    INIT_05 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
    INIT_06 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
    INIT_07 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
    INIT_08 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
    INIT_09 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
    INIT_0A : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
    INIT_0B : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
    INIT_0C : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
    INIT_0D : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
    INIT_0E : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
    INIT_0F : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
    INIT_10 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
    INIT_11 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
    INIT_12 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
    INIT_13 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
    INIT_14 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
    INIT_15 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
    INIT_16 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
    INIT_17 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
    INIT_18 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
    INIT_19 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
    INIT_1A : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
    INIT_1B : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
    INIT_1C : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
    INIT_1D : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
    INIT_1E : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
    INIT_1F : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
    INIT_20 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
    INIT_21 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
    INIT_22 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
    INIT_23 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
    INIT_24 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
    INIT_25 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
    INIT_26 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
    INIT_27 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
    INIT_28 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
    INIT_29 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
    INIT_2A : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
    INIT_2B : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
    INIT_2C : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
    INIT_2D : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
    INIT_2E : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
    INIT_2F : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
    INIT_30 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
    INIT_31 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
    INIT_32 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
    INIT_33 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
    INIT_34 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
    INIT_35 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
    INIT_36 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
    INIT_37 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
    INIT_38 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
    INIT_39 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
    INIT_3A : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
    INIT_3B : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
    INIT_3C : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
    INIT_3D : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
    INIT_3E : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
    INIT_3F : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000" );
  PORT (
    DO : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    DOP : OUT STD_LOGIC_VECTOR (0 DOWNTO 0);    
    DI : IN STD_LOGIC_VECTOR (7 DOWNTO 0); 
    DIP : IN STD_LOGIC_VECTOR (0 DOWNTO 0);     
    ADDR : IN STD_LOGIC_VECTOR (10 DOWNTO 0);
    CLK : IN STD_ULOGIC;
    EN : IN STD_ULOGIC;
    SSR : IN STD_ULOGIC;
    WE : IN STD_ULOGIC ); 
  END COMPONENT;  

  COMPONENT pulse 
  PORT (
    clk: IN STD_LOGIC;
    clr: IN STD_LOGIC;
    pulse_i: IN STD_LOGIC;
    pulse_o: OUT STD_LOGIC;
    pulse_d: OUT STD_LOGIC );
  END COMPONENT;  
  
  SIGNAL rom_bram_00_dat_o : STD_LOGIC_VECTOR (7 DOWNTO 0); 
  SIGNAL rom_bram_01_dat_o : STD_LOGIC_VECTOR (7 DOWNTO 0); 
  SIGNAL rom_bram_02_dat_o : STD_LOGIC_VECTOR (7 DOWNTO 0); 
  SIGNAL rom_bram_03_dat_o : STD_LOGIC_VECTOR (7 DOWNTO 0); 
  SIGNAL rom_bram_04_dat_o : STD_LOGIC_VECTOR (7 DOWNTO 0); 
  SIGNAL rom_bram_05_dat_o : STD_LOGIC_VECTOR (7 DOWNTO 0); 
  SIGNAL rom_bram_06_dat_o : STD_LOGIC_VECTOR (7 DOWNTO 0); 
  SIGNAL rom_bram_07_dat_o : STD_LOGIC_VECTOR (7 DOWNTO 0); 
  SIGNAL rom_bram_08_dat_o : STD_LOGIC_VECTOR (7 DOWNTO 0); 
  SIGNAL rom_bram_09_dat_o : STD_LOGIC_VECTOR (7 DOWNTO 0); 
  SIGNAL rom_bram_0A_dat_o : STD_LOGIC_VECTOR (7 DOWNTO 0); 
  SIGNAL rom_bram_0B_dat_o : STD_LOGIC_VECTOR (7 DOWNTO 0); 
  SIGNAL rom_bram_0C_dat_o : STD_LOGIC_VECTOR (7 DOWNTO 0); 
  SIGNAL rom_bram_0D_dat_o : STD_LOGIC_VECTOR (7 DOWNTO 0); 
  SIGNAL rom_bram_0E_dat_o : STD_LOGIC_VECTOR (7 DOWNTO 0); 
  SIGNAL rom_bram_0F_dat_o : STD_LOGIC_VECTOR (7 DOWNTO 0); 
  SIGNAL rom_bram_10_dat_o : STD_LOGIC_VECTOR (7 DOWNTO 0); 
  SIGNAL rom_bram_11_dat_o : STD_LOGIC_VECTOR (7 DOWNTO 0); 
  SIGNAL rom_bram_12_dat_o : STD_LOGIC_VECTOR (7 DOWNTO 0); 
  SIGNAL rom_bram_13_dat_o : STD_LOGIC_VECTOR (7 DOWNTO 0); 
  SIGNAL rom_bram_14_dat_o : STD_LOGIC_VECTOR (7 DOWNTO 0); 
  SIGNAL rom_bram_15_dat_o : STD_LOGIC_VECTOR (7 DOWNTO 0); 
  SIGNAL rom_bram_16_dat_o : STD_LOGIC_VECTOR (7 DOWNTO 0); 
  SIGNAL rom_bram_17_dat_o : STD_LOGIC_VECTOR (7 DOWNTO 0); 
  SIGNAL rom_bram_18_dat_o : STD_LOGIC_VECTOR (7 DOWNTO 0); 
  SIGNAL rom_bram_19_dat_o : STD_LOGIC_VECTOR (7 DOWNTO 0); 
  SIGNAL rom_bram_1A_dat_o : STD_LOGIC_VECTOR (7 DOWNTO 0); 
  SIGNAL rom_bram_1B_dat_o : STD_LOGIC_VECTOR (7 DOWNTO 0); 
  SIGNAL rom_bram_1C_dat_o : STD_LOGIC_VECTOR (7 DOWNTO 0); 
  SIGNAL rom_bram_1D_dat_o : STD_LOGIC_VECTOR (7 DOWNTO 0); 
  SIGNAL rom_bram_1E_dat_o : STD_LOGIC_VECTOR (7 DOWNTO 0); 
  SIGNAL rom_bram_1F_dat_o : STD_LOGIC_VECTOR (7 DOWNTO 0);
  
  SIGNAL ack_int : STD_LOGIC;

BEGIN

  --
  -- signal buffers
  --
  
  ack_int <= stb_i and cyc_i and not rst_i;

  --
  -- processes
  --

  mux : PROCESS (adr_i,
                 rom_bram_00_dat_o, rom_bram_01_dat_o, rom_bram_02_dat_o, rom_bram_03_dat_o,
                 rom_bram_04_dat_o, rom_bram_05_dat_o, rom_bram_06_dat_o, rom_bram_07_dat_o,  
                 rom_bram_08_dat_o, rom_bram_09_dat_o, rom_bram_0A_dat_o, rom_bram_0B_dat_o, 
                 rom_bram_0C_dat_o, rom_bram_0D_dat_o, rom_bram_0E_dat_o, rom_bram_0F_dat_o, 
                 rom_bram_10_dat_o, rom_bram_11_dat_o, rom_bram_12_dat_o, rom_bram_13_dat_o,  
                 rom_bram_14_dat_o, rom_bram_15_dat_o, rom_bram_16_dat_o, rom_bram_17_dat_o, 
                 rom_bram_18_dat_o, rom_bram_19_dat_o, rom_bram_1A_dat_o, rom_bram_1B_dat_o, 
                 rom_bram_1C_dat_o, rom_bram_1D_dat_o, rom_bram_1E_dat_o, rom_bram_1F_dat_o )
  BEGIN
    CASE adr_i(15 DOWNTO 11) is
      WHEN "00000" => dat_o <= rom_bram_00_dat_o;
      WHEN "00001" => dat_o <= rom_bram_01_dat_o;
      WHEN "00010" => dat_o <= rom_bram_02_dat_o;
      WHEN "00011" => dat_o <= rom_bram_03_dat_o;
      WHEN "00100" => dat_o <= rom_bram_04_dat_o;
      WHEN "00101" => dat_o <= rom_bram_05_dat_o;
      WHEN "00110" => dat_o <= rom_bram_06_dat_o;
      WHEN "00111" => dat_o <= rom_bram_07_dat_o;
      WHEN "01000" => dat_o <= rom_bram_08_dat_o;
      WHEN "01001" => dat_o <= rom_bram_09_dat_o;
      WHEN "01010" => dat_o <= rom_bram_0A_dat_o;
      WHEN "01011" => dat_o <= rom_bram_0B_dat_o;
      WHEN "01100" => dat_o <= rom_bram_0C_dat_o;
      WHEN "01101" => dat_o <= rom_bram_0D_dat_o;
      WHEN "01110" => dat_o <= rom_bram_0E_dat_o;
      WHEN "01111" => dat_o <= rom_bram_0F_dat_o;
      WHEN "10000" => dat_o <= rom_bram_10_dat_o;
      WHEN "10001" => dat_o <= rom_bram_11_dat_o;
      WHEN "10010" => dat_o <= rom_bram_12_dat_o;
      WHEN "10011" => dat_o <= rom_bram_13_dat_o;
      WHEN "10100" => dat_o <= rom_bram_14_dat_o;
      WHEN "10101" => dat_o <= rom_bram_15_dat_o;
      WHEN "10110" => dat_o <= rom_bram_16_dat_o;
      WHEN "10111" => dat_o <= rom_bram_17_dat_o;
      WHEN "11000" => dat_o <= rom_bram_18_dat_o;
      WHEN "11001" => dat_o <= rom_bram_19_dat_o;
      WHEN "11010" => dat_o <= rom_bram_1A_dat_o;
      WHEN "11011" => dat_o <= rom_bram_1B_dat_o;
      WHEN "11100" => dat_o <= rom_bram_1C_dat_o;
      WHEN "11101" => dat_o <= rom_bram_1D_dat_o;
      WHEN "11110" => dat_o <= rom_bram_1E_dat_o;
      WHEN "11111" => dat_o <= rom_bram_1F_dat_o;
      WHEN OTHERS  => dat_o <= (OTHERS=>'0');
    END CASE;
  END PROCESS;       
  --
  -- components
  --

  ack_pulse : pulse PORT MAP(
    clk => clk_i,
    clr => rst_i,
    pulse_i => ack_int,
    pulse_o => ack_o,
    pulse_d => OPEN );
    
  
  -- BRAM 0 in address space [0x00000000:0x000007FF], bit lane [7:0]
  rom_bram_00 : RAMB16_S9 
  GENERIC MAP(
    INIT_00 => rom_bram_00_INIT_00,
    INIT_01 => rom_bram_00_INIT_01,
    INIT_02 => rom_bram_00_INIT_02,
    INIT_03 => rom_bram_00_INIT_03,
    INIT_04 => rom_bram_00_INIT_04,
    INIT_05 => rom_bram_00_INIT_05,
    INIT_06 => rom_bram_00_INIT_06,
    INIT_07 => rom_bram_00_INIT_07,
    INIT_08 => rom_bram_00_INIT_08,
    INIT_09 => rom_bram_00_INIT_09,
    INIT_0A => rom_bram_00_INIT_0A,
    INIT_0B => rom_bram_00_INIT_0B,
    INIT_0C => rom_bram_00_INIT_0C,
    INIT_0D => rom_bram_00_INIT_0D,
    INIT_0E => rom_bram_00_INIT_0E,
    INIT_0F => rom_bram_00_INIT_0F,
    INIT_10 => rom_bram_00_INIT_10,
    INIT_11 => rom_bram_00_INIT_11,
    INIT_12 => rom_bram_00_INIT_12,
    INIT_13 => rom_bram_00_INIT_13,
    INIT_14 => rom_bram_00_INIT_14,
    INIT_15 => rom_bram_00_INIT_15,
    INIT_16 => rom_bram_00_INIT_16,
    INIT_17 => rom_bram_00_INIT_17,
    INIT_18 => rom_bram_00_INIT_18,
    INIT_19 => rom_bram_00_INIT_19,
    INIT_1A => rom_bram_00_INIT_1A,
    INIT_1B => rom_bram_00_INIT_1B,
    INIT_1C => rom_bram_00_INIT_1C,
    INIT_1D => rom_bram_00_INIT_1D,
    INIT_1E => rom_bram_00_INIT_1E,
    INIT_1F => rom_bram_00_INIT_1F,
    INIT_20 => rom_bram_00_INIT_20,
    INIT_21 => rom_bram_00_INIT_21,
    INIT_22 => rom_bram_00_INIT_22,
    INIT_23 => rom_bram_00_INIT_23,
    INIT_24 => rom_bram_00_INIT_24,
    INIT_25 => rom_bram_00_INIT_25,
    INIT_26 => rom_bram_00_INIT_26,
    INIT_27 => rom_bram_00_INIT_27,
    INIT_28 => rom_bram_00_INIT_28,
    INIT_29 => rom_bram_00_INIT_29,
    INIT_2A => rom_bram_00_INIT_2A,
    INIT_2B => rom_bram_00_INIT_2B,
    INIT_2C => rom_bram_00_INIT_2C,
    INIT_2D => rom_bram_00_INIT_2D,
    INIT_2E => rom_bram_00_INIT_2E,
    INIT_2F => rom_bram_00_INIT_2F,
    INIT_30 => rom_bram_00_INIT_30,
    INIT_31 => rom_bram_00_INIT_31,
    INIT_32 => rom_bram_00_INIT_32,
    INIT_33 => rom_bram_00_INIT_33,
    INIT_34 => rom_bram_00_INIT_34,
    INIT_35 => rom_bram_00_INIT_35,
    INIT_36 => rom_bram_00_INIT_36,
    INIT_37 => rom_bram_00_INIT_37,
    INIT_38 => rom_bram_00_INIT_38,
    INIT_39 => rom_bram_00_INIT_39,
    INIT_3A => rom_bram_00_INIT_3A,
    INIT_3B => rom_bram_00_INIT_3B,
    INIT_3C => rom_bram_00_INIT_3C,
    INIT_3D => rom_bram_00_INIT_3D,
    INIT_3E => rom_bram_00_INIT_3E,
    INIT_3F => rom_bram_00_INIT_3F )
  PORT MAP( 
    DO => rom_bram_00_dat_o,
    dop => OPEN,    
    di => "00000000",
    dip => "0",
    addr => adr_i(10 DOWNTO 0), 
    clk => clk_i,    
    en => '1',
    ssr => '0',
    we => '0' );

  -- BRAM 1 in address space [0x00000800:0x00000FFF], bit lane [7:0]
  rom_bram_01 : RAMB16_S9 
  GENERIC MAP(
    INIT_00 => rom_bram_01_INIT_00,
    INIT_01 => rom_bram_01_INIT_01,
    INIT_02 => rom_bram_01_INIT_02,
    INIT_03 => rom_bram_01_INIT_03,
    INIT_04 => rom_bram_01_INIT_04,
    INIT_05 => rom_bram_01_INIT_05,
    INIT_06 => rom_bram_01_INIT_06,
    INIT_07 => rom_bram_01_INIT_07,
    INIT_08 => rom_bram_01_INIT_08,
    INIT_09 => rom_bram_01_INIT_09,
    INIT_0A => rom_bram_01_INIT_0A,
    INIT_0B => rom_bram_01_INIT_0B,
    INIT_0C => rom_bram_01_INIT_0C,
    INIT_0D => rom_bram_01_INIT_0D,
    INIT_0E => rom_bram_01_INIT_0E,
    INIT_0F => rom_bram_01_INIT_0F,
    INIT_10 => rom_bram_01_INIT_10,
    INIT_11 => rom_bram_01_INIT_11,
    INIT_12 => rom_bram_01_INIT_12,
    INIT_13 => rom_bram_01_INIT_13,
    INIT_14 => rom_bram_01_INIT_14,
    INIT_15 => rom_bram_01_INIT_15,
    INIT_16 => rom_bram_01_INIT_16,
    INIT_17 => rom_bram_01_INIT_17,
    INIT_18 => rom_bram_01_INIT_18,
    INIT_19 => rom_bram_01_INIT_19,
    INIT_1A => rom_bram_01_INIT_1A,
    INIT_1B => rom_bram_01_INIT_1B,
    INIT_1C => rom_bram_01_INIT_1C,
    INIT_1D => rom_bram_01_INIT_1D,
    INIT_1E => rom_bram_01_INIT_1E,
    INIT_1F => rom_bram_01_INIT_1F,
    INIT_20 => rom_bram_01_INIT_20,
    INIT_21 => rom_bram_01_INIT_21,
    INIT_22 => rom_bram_01_INIT_22,
    INIT_23 => rom_bram_01_INIT_23,
    INIT_24 => rom_bram_01_INIT_24,
    INIT_25 => rom_bram_01_INIT_25,
    INIT_26 => rom_bram_01_INIT_26,
    INIT_27 => rom_bram_01_INIT_27,
    INIT_28 => rom_bram_01_INIT_28,
    INIT_29 => rom_bram_01_INIT_29,
    INIT_2A => rom_bram_01_INIT_2A,
    INIT_2B => rom_bram_01_INIT_2B,
    INIT_2C => rom_bram_01_INIT_2C,
    INIT_2D => rom_bram_01_INIT_2D,
    INIT_2E => rom_bram_01_INIT_2E,
    INIT_2F => rom_bram_01_INIT_2F,
    INIT_30 => rom_bram_01_INIT_30,
    INIT_31 => rom_bram_01_INIT_31,
    INIT_32 => rom_bram_01_INIT_32,
    INIT_33 => rom_bram_01_INIT_33,
    INIT_34 => rom_bram_01_INIT_34,
    INIT_35 => rom_bram_01_INIT_35,
    INIT_36 => rom_bram_01_INIT_36,
    INIT_37 => rom_bram_01_INIT_37,
    INIT_38 => rom_bram_01_INIT_38,
    INIT_39 => rom_bram_01_INIT_39,
    INIT_3A => rom_bram_01_INIT_3A,
    INIT_3B => rom_bram_01_INIT_3B,
    INIT_3C => rom_bram_01_INIT_3C,
    INIT_3D => rom_bram_01_INIT_3D,
    INIT_3E => rom_bram_01_INIT_3E,
    INIT_3F => rom_bram_01_INIT_3F )
  PORT MAP( 
    DO => rom_bram_01_dat_o,
    dop => OPEN,    
    di => "00000000",
    dip => "0",
    addr => adr_i(10 DOWNTO 0), 
    clk => clk_i,    
    en => '1',
    ssr => '0',
    we => '0' );
    
  -- BRAM 2 in address space [0x00001000:0x000017FF], bit lane [7:0]
  rom_bram_02 : RAMB16_S9 
  GENERIC MAP(
    INIT_00 => rom_bram_02_INIT_00,
    INIT_01 => rom_bram_02_INIT_01,
    INIT_02 => rom_bram_02_INIT_02,
    INIT_03 => rom_bram_02_INIT_03,
    INIT_04 => rom_bram_02_INIT_04,
    INIT_05 => rom_bram_02_INIT_05,
    INIT_06 => rom_bram_02_INIT_06,
    INIT_07 => rom_bram_02_INIT_07,
    INIT_08 => rom_bram_02_INIT_08,
    INIT_09 => rom_bram_02_INIT_09,
    INIT_0A => rom_bram_02_INIT_0A,
    INIT_0B => rom_bram_02_INIT_0B,
    INIT_0C => rom_bram_02_INIT_0C,
    INIT_0D => rom_bram_02_INIT_0D,
    INIT_0E => rom_bram_02_INIT_0E,
    INIT_0F => rom_bram_02_INIT_0F,
    INIT_10 => rom_bram_02_INIT_10,
    INIT_11 => rom_bram_02_INIT_11,
    INIT_12 => rom_bram_02_INIT_12,
    INIT_13 => rom_bram_02_INIT_13,
    INIT_14 => rom_bram_02_INIT_14,
    INIT_15 => rom_bram_02_INIT_15,
    INIT_16 => rom_bram_02_INIT_16,
    INIT_17 => rom_bram_02_INIT_17,
    INIT_18 => rom_bram_02_INIT_18,
    INIT_19 => rom_bram_02_INIT_19,
    INIT_1A => rom_bram_02_INIT_1A,
    INIT_1B => rom_bram_02_INIT_1B,
    INIT_1C => rom_bram_02_INIT_1C,
    INIT_1D => rom_bram_02_INIT_1D,
    INIT_1E => rom_bram_02_INIT_1E,
    INIT_1F => rom_bram_02_INIT_1F,
    INIT_20 => rom_bram_02_INIT_20,
    INIT_21 => rom_bram_02_INIT_21,
    INIT_22 => rom_bram_02_INIT_22,
    INIT_23 => rom_bram_02_INIT_23,
    INIT_24 => rom_bram_02_INIT_24,
    INIT_25 => rom_bram_02_INIT_25,
    INIT_26 => rom_bram_02_INIT_26,
    INIT_27 => rom_bram_02_INIT_27,
    INIT_28 => rom_bram_02_INIT_28,
    INIT_29 => rom_bram_02_INIT_29,
    INIT_2A => rom_bram_02_INIT_2A,
    INIT_2B => rom_bram_02_INIT_2B,
    INIT_2C => rom_bram_02_INIT_2C,
    INIT_2D => rom_bram_02_INIT_2D,
    INIT_2E => rom_bram_02_INIT_2E,
    INIT_2F => rom_bram_02_INIT_2F,
    INIT_30 => rom_bram_02_INIT_30,
    INIT_31 => rom_bram_02_INIT_31,
    INIT_32 => rom_bram_02_INIT_32,
    INIT_33 => rom_bram_02_INIT_33,
    INIT_34 => rom_bram_02_INIT_34,
    INIT_35 => rom_bram_02_INIT_35,
    INIT_36 => rom_bram_02_INIT_36,
    INIT_37 => rom_bram_02_INIT_37,
    INIT_38 => rom_bram_02_INIT_38,
    INIT_39 => rom_bram_02_INIT_39,
    INIT_3A => rom_bram_02_INIT_3A,
    INIT_3B => rom_bram_02_INIT_3B,
    INIT_3C => rom_bram_02_INIT_3C,
    INIT_3D => rom_bram_02_INIT_3D,
    INIT_3E => rom_bram_02_INIT_3E,
    INIT_3F => rom_bram_02_INIT_3F )
  PORT MAP( 
    DO => rom_bram_02_dat_o,
    dop => OPEN,    
    di => "00000000",
    dip => "0",
    addr => adr_i(10 DOWNTO 0), 
    clk => clk_i,    
    en => '1',
    ssr => '0',
    we => '0' );
    
  -- BRAM 3 in address space [0x00001800:0x00001FFF], bit lane [7:0]
  rom_bram_03 : RAMB16_S9 
  GENERIC MAP(
    INIT_00 => rom_bram_03_INIT_00,
    INIT_01 => rom_bram_03_INIT_01,
    INIT_02 => rom_bram_03_INIT_02,
    INIT_03 => rom_bram_03_INIT_03,
    INIT_04 => rom_bram_03_INIT_04,
    INIT_05 => rom_bram_03_INIT_05,
    INIT_06 => rom_bram_03_INIT_06,
    INIT_07 => rom_bram_03_INIT_07,
    INIT_08 => rom_bram_03_INIT_08,
    INIT_09 => rom_bram_03_INIT_09,
    INIT_0A => rom_bram_03_INIT_0A,
    INIT_0B => rom_bram_03_INIT_0B,
    INIT_0C => rom_bram_03_INIT_0C,
    INIT_0D => rom_bram_03_INIT_0D,
    INIT_0E => rom_bram_03_INIT_0E,
    INIT_0F => rom_bram_03_INIT_0F,
    INIT_10 => rom_bram_03_INIT_10,
    INIT_11 => rom_bram_03_INIT_11,
    INIT_12 => rom_bram_03_INIT_12,
    INIT_13 => rom_bram_03_INIT_13,
    INIT_14 => rom_bram_03_INIT_14,
    INIT_15 => rom_bram_03_INIT_15,
    INIT_16 => rom_bram_03_INIT_16,
    INIT_17 => rom_bram_03_INIT_17,
    INIT_18 => rom_bram_03_INIT_18,
    INIT_19 => rom_bram_03_INIT_19,
    INIT_1A => rom_bram_03_INIT_1A,
    INIT_1B => rom_bram_03_INIT_1B,
    INIT_1C => rom_bram_03_INIT_1C,
    INIT_1D => rom_bram_03_INIT_1D,
    INIT_1E => rom_bram_03_INIT_1E,
    INIT_1F => rom_bram_03_INIT_1F,
    INIT_20 => rom_bram_03_INIT_20,
    INIT_21 => rom_bram_03_INIT_21,
    INIT_22 => rom_bram_03_INIT_22,
    INIT_23 => rom_bram_03_INIT_23,
    INIT_24 => rom_bram_03_INIT_24,
    INIT_25 => rom_bram_03_INIT_25,
    INIT_26 => rom_bram_03_INIT_26,
    INIT_27 => rom_bram_03_INIT_27,
    INIT_28 => rom_bram_03_INIT_28,
    INIT_29 => rom_bram_03_INIT_29,
    INIT_2A => rom_bram_03_INIT_2A,
    INIT_2B => rom_bram_03_INIT_2B,
    INIT_2C => rom_bram_03_INIT_2C,
    INIT_2D => rom_bram_03_INIT_2D,
    INIT_2E => rom_bram_03_INIT_2E,
    INIT_2F => rom_bram_03_INIT_2F,
    INIT_30 => rom_bram_03_INIT_30,
    INIT_31 => rom_bram_03_INIT_31,
    INIT_32 => rom_bram_03_INIT_32,
    INIT_33 => rom_bram_03_INIT_33,
    INIT_34 => rom_bram_03_INIT_34,
    INIT_35 => rom_bram_03_INIT_35,
    INIT_36 => rom_bram_03_INIT_36,
    INIT_37 => rom_bram_03_INIT_37,
    INIT_38 => rom_bram_03_INIT_38,
    INIT_39 => rom_bram_03_INIT_39,
    INIT_3A => rom_bram_03_INIT_3A,
    INIT_3B => rom_bram_03_INIT_3B,
    INIT_3C => rom_bram_03_INIT_3C,
    INIT_3D => rom_bram_03_INIT_3D,
    INIT_3E => rom_bram_03_INIT_3E,
    INIT_3F => rom_bram_03_INIT_3F )
  PORT MAP( 
    DO => rom_bram_03_dat_o,
    dop => OPEN,    
    di => "00000000",
    dip => "0",
    addr => adr_i(10 DOWNTO 0), 
    clk => clk_i,    
    en => '1',
    ssr => '0',
    we => '0' ); 
  
  -- BRAM 4 in address space [0x00002000:0x000027FF], bit lane [7:0]
  rom_bram_04 : RAMB16_S9 
  GENERIC MAP(
    INIT_00 => rom_bram_04_INIT_00,
    INIT_01 => rom_bram_04_INIT_01,
    INIT_02 => rom_bram_04_INIT_02,
    INIT_03 => rom_bram_04_INIT_03,
    INIT_04 => rom_bram_04_INIT_04,
    INIT_05 => rom_bram_04_INIT_05,
    INIT_06 => rom_bram_04_INIT_06,
    INIT_07 => rom_bram_04_INIT_07,
    INIT_08 => rom_bram_04_INIT_08,
    INIT_09 => rom_bram_04_INIT_09,
    INIT_0A => rom_bram_04_INIT_0A,
    INIT_0B => rom_bram_04_INIT_0B,
    INIT_0C => rom_bram_04_INIT_0C,
    INIT_0D => rom_bram_04_INIT_0D,
    INIT_0E => rom_bram_04_INIT_0E,
    INIT_0F => rom_bram_04_INIT_0F,
    INIT_10 => rom_bram_04_INIT_10,
    INIT_11 => rom_bram_04_INIT_11,
    INIT_12 => rom_bram_04_INIT_12,
    INIT_13 => rom_bram_04_INIT_13,
    INIT_14 => rom_bram_04_INIT_14,
    INIT_15 => rom_bram_04_INIT_15,
    INIT_16 => rom_bram_04_INIT_16,
    INIT_17 => rom_bram_04_INIT_17,
    INIT_18 => rom_bram_04_INIT_18,
    INIT_19 => rom_bram_04_INIT_19,
    INIT_1A => rom_bram_04_INIT_1A,
    INIT_1B => rom_bram_04_INIT_1B,
    INIT_1C => rom_bram_04_INIT_1C,
    INIT_1D => rom_bram_04_INIT_1D,
    INIT_1E => rom_bram_04_INIT_1E,
    INIT_1F => rom_bram_04_INIT_1F,
    INIT_20 => rom_bram_04_INIT_20,
    INIT_21 => rom_bram_04_INIT_21,
    INIT_22 => rom_bram_04_INIT_22,
    INIT_23 => rom_bram_04_INIT_23,
    INIT_24 => rom_bram_04_INIT_24,
    INIT_25 => rom_bram_04_INIT_25,
    INIT_26 => rom_bram_04_INIT_26,
    INIT_27 => rom_bram_04_INIT_27,
    INIT_28 => rom_bram_04_INIT_28,
    INIT_29 => rom_bram_04_INIT_29,
    INIT_2A => rom_bram_04_INIT_2A,
    INIT_2B => rom_bram_04_INIT_2B,
    INIT_2C => rom_bram_04_INIT_2C,
    INIT_2D => rom_bram_04_INIT_2D,
    INIT_2E => rom_bram_04_INIT_2E,
    INIT_2F => rom_bram_04_INIT_2F,
    INIT_30 => rom_bram_04_INIT_30,
    INIT_31 => rom_bram_04_INIT_31,
    INIT_32 => rom_bram_04_INIT_32,
    INIT_33 => rom_bram_04_INIT_33,
    INIT_34 => rom_bram_04_INIT_34,
    INIT_35 => rom_bram_04_INIT_35,
    INIT_36 => rom_bram_04_INIT_36,
    INIT_37 => rom_bram_04_INIT_37,
    INIT_38 => rom_bram_04_INIT_38,
    INIT_39 => rom_bram_04_INIT_39,
    INIT_3A => rom_bram_04_INIT_3A,
    INIT_3B => rom_bram_04_INIT_3B,
    INIT_3C => rom_bram_04_INIT_3C,
    INIT_3D => rom_bram_04_INIT_3D,
    INIT_3E => rom_bram_04_INIT_3E,
    INIT_3F => rom_bram_04_INIT_3F )
  PORT MAP( 
    DO => rom_bram_04_dat_o,
    dop => OPEN,    
    di => "00000000",
    dip => "0",
    addr => adr_i(10 DOWNTO 0), 
    clk => clk_i,    
    en => '1',
    ssr => '0',
    we => '0' );

  -- BRAM 5 in address space [0x00002800:0x00002FFF], bit lane [7:0]
  rom_bram_05 : RAMB16_S9 
  GENERIC MAP(
    INIT_00 => rom_bram_05_INIT_00,
    INIT_01 => rom_bram_05_INIT_01,
    INIT_02 => rom_bram_05_INIT_02,
    INIT_03 => rom_bram_05_INIT_03,
    INIT_04 => rom_bram_05_INIT_04,
    INIT_05 => rom_bram_05_INIT_05,
    INIT_06 => rom_bram_05_INIT_06,
    INIT_07 => rom_bram_05_INIT_07,
    INIT_08 => rom_bram_05_INIT_08,
    INIT_09 => rom_bram_05_INIT_09,
    INIT_0A => rom_bram_05_INIT_0A,
    INIT_0B => rom_bram_05_INIT_0B,
    INIT_0C => rom_bram_05_INIT_0C,
    INIT_0D => rom_bram_05_INIT_0D,
    INIT_0E => rom_bram_05_INIT_0E,
    INIT_0F => rom_bram_05_INIT_0F,
    INIT_10 => rom_bram_05_INIT_10,
    INIT_11 => rom_bram_05_INIT_11,
    INIT_12 => rom_bram_05_INIT_12,
    INIT_13 => rom_bram_05_INIT_13,
    INIT_14 => rom_bram_05_INIT_14,
    INIT_15 => rom_bram_05_INIT_15,
    INIT_16 => rom_bram_05_INIT_16,
    INIT_17 => rom_bram_05_INIT_17,
    INIT_18 => rom_bram_05_INIT_18,
    INIT_19 => rom_bram_05_INIT_19,
    INIT_1A => rom_bram_05_INIT_1A,
    INIT_1B => rom_bram_05_INIT_1B,
    INIT_1C => rom_bram_05_INIT_1C,
    INIT_1D => rom_bram_05_INIT_1D,
    INIT_1E => rom_bram_05_INIT_1E,
    INIT_1F => rom_bram_05_INIT_1F,
    INIT_20 => rom_bram_05_INIT_20,
    INIT_21 => rom_bram_05_INIT_21,
    INIT_22 => rom_bram_05_INIT_22,
    INIT_23 => rom_bram_05_INIT_23,
    INIT_24 => rom_bram_05_INIT_24,
    INIT_25 => rom_bram_05_INIT_25,
    INIT_26 => rom_bram_05_INIT_26,
    INIT_27 => rom_bram_05_INIT_27,
    INIT_28 => rom_bram_05_INIT_28,
    INIT_29 => rom_bram_05_INIT_29,
    INIT_2A => rom_bram_05_INIT_2A,
    INIT_2B => rom_bram_05_INIT_2B,
    INIT_2C => rom_bram_05_INIT_2C,
    INIT_2D => rom_bram_05_INIT_2D,
    INIT_2E => rom_bram_05_INIT_2E,
    INIT_2F => rom_bram_05_INIT_2F,
    INIT_30 => rom_bram_05_INIT_30,
    INIT_31 => rom_bram_05_INIT_31,
    INIT_32 => rom_bram_05_INIT_32,
    INIT_33 => rom_bram_05_INIT_33,
    INIT_34 => rom_bram_05_INIT_34,
    INIT_35 => rom_bram_05_INIT_35,
    INIT_36 => rom_bram_05_INIT_36,
    INIT_37 => rom_bram_05_INIT_37,
    INIT_38 => rom_bram_05_INIT_38,
    INIT_39 => rom_bram_05_INIT_39,
    INIT_3A => rom_bram_05_INIT_3A,
    INIT_3B => rom_bram_05_INIT_3B,
    INIT_3C => rom_bram_05_INIT_3C,
    INIT_3D => rom_bram_05_INIT_3D,
    INIT_3E => rom_bram_05_INIT_3E,
    INIT_3F => rom_bram_05_INIT_3F )
  PORT MAP( 
    DO => rom_bram_05_dat_o,
    dop => OPEN,    
    di => "00000000",
    dip => "0",
    addr => adr_i(10 DOWNTO 0), 
    clk => clk_i,    
    en => '1',
    ssr => '0',
    we => '0' );
    
  -- BRAM 6 in address space [0x00003000:0x000037FF], bit lane [7:0]
  rom_bram_06 : RAMB16_S9 
  GENERIC MAP(
    INIT_00 => rom_bram_06_INIT_00,
    INIT_01 => rom_bram_06_INIT_01,
    INIT_02 => rom_bram_06_INIT_02,
    INIT_03 => rom_bram_06_INIT_03,
    INIT_04 => rom_bram_06_INIT_04,
    INIT_05 => rom_bram_06_INIT_05,
    INIT_06 => rom_bram_06_INIT_06,
    INIT_07 => rom_bram_06_INIT_07,
    INIT_08 => rom_bram_06_INIT_08,
    INIT_09 => rom_bram_06_INIT_09,
    INIT_0A => rom_bram_06_INIT_0A,
    INIT_0B => rom_bram_06_INIT_0B,
    INIT_0C => rom_bram_06_INIT_0C,
    INIT_0D => rom_bram_06_INIT_0D,
    INIT_0E => rom_bram_06_INIT_0E,
    INIT_0F => rom_bram_06_INIT_0F,
    INIT_10 => rom_bram_06_INIT_10,
    INIT_11 => rom_bram_06_INIT_11,
    INIT_12 => rom_bram_06_INIT_12,
    INIT_13 => rom_bram_06_INIT_13,
    INIT_14 => rom_bram_06_INIT_14,
    INIT_15 => rom_bram_06_INIT_15,
    INIT_16 => rom_bram_06_INIT_16,
    INIT_17 => rom_bram_06_INIT_17,
    INIT_18 => rom_bram_06_INIT_18,
    INIT_19 => rom_bram_06_INIT_19,
    INIT_1A => rom_bram_06_INIT_1A,
    INIT_1B => rom_bram_06_INIT_1B,
    INIT_1C => rom_bram_06_INIT_1C,
    INIT_1D => rom_bram_06_INIT_1D,
    INIT_1E => rom_bram_06_INIT_1E,
    INIT_1F => rom_bram_06_INIT_1F,
    INIT_20 => rom_bram_06_INIT_20,
    INIT_21 => rom_bram_06_INIT_21,
    INIT_22 => rom_bram_06_INIT_22,
    INIT_23 => rom_bram_06_INIT_23,
    INIT_24 => rom_bram_06_INIT_24,
    INIT_25 => rom_bram_06_INIT_25,
    INIT_26 => rom_bram_06_INIT_26,
    INIT_27 => rom_bram_06_INIT_27,
    INIT_28 => rom_bram_06_INIT_28,
    INIT_29 => rom_bram_06_INIT_29,
    INIT_2A => rom_bram_06_INIT_2A,
    INIT_2B => rom_bram_06_INIT_2B,
    INIT_2C => rom_bram_06_INIT_2C,
    INIT_2D => rom_bram_06_INIT_2D,
    INIT_2E => rom_bram_06_INIT_2E,
    INIT_2F => rom_bram_06_INIT_2F,
    INIT_30 => rom_bram_06_INIT_30,
    INIT_31 => rom_bram_06_INIT_31,
    INIT_32 => rom_bram_06_INIT_32,
    INIT_33 => rom_bram_06_INIT_33,
    INIT_34 => rom_bram_06_INIT_34,
    INIT_35 => rom_bram_06_INIT_35,
    INIT_36 => rom_bram_06_INIT_36,
    INIT_37 => rom_bram_06_INIT_37,
    INIT_38 => rom_bram_06_INIT_38,
    INIT_39 => rom_bram_06_INIT_39,
    INIT_3A => rom_bram_06_INIT_3A,
    INIT_3B => rom_bram_06_INIT_3B,
    INIT_3C => rom_bram_06_INIT_3C,
    INIT_3D => rom_bram_06_INIT_3D,
    INIT_3E => rom_bram_06_INIT_3E,
    INIT_3F => rom_bram_06_INIT_3F )
  PORT MAP( 
    DO => rom_bram_06_dat_o,
    dop => OPEN,    
    di => "00000000",
    dip => "0",
    addr => adr_i(10 DOWNTO 0), 
    clk => clk_i,    
    en => '1',
    ssr => '0',
    we => '0' );
    
  -- BRAM 7 in address space [0x00003800:0x00003FFF], bit lane [7:0]
  rom_bram_07 : RAMB16_S9 
  GENERIC MAP(
    INIT_00 => rom_bram_07_INIT_00,
    INIT_01 => rom_bram_07_INIT_01,
    INIT_02 => rom_bram_07_INIT_02,
    INIT_03 => rom_bram_07_INIT_03,
    INIT_04 => rom_bram_07_INIT_04,
    INIT_05 => rom_bram_07_INIT_05,
    INIT_06 => rom_bram_07_INIT_06,
    INIT_07 => rom_bram_07_INIT_07,
    INIT_08 => rom_bram_07_INIT_08,
    INIT_09 => rom_bram_07_INIT_09,
    INIT_0A => rom_bram_07_INIT_0A,
    INIT_0B => rom_bram_07_INIT_0B,
    INIT_0C => rom_bram_07_INIT_0C,
    INIT_0D => rom_bram_07_INIT_0D,
    INIT_0E => rom_bram_07_INIT_0E,
    INIT_0F => rom_bram_07_INIT_0F,
    INIT_10 => rom_bram_07_INIT_10,
    INIT_11 => rom_bram_07_INIT_11,
    INIT_12 => rom_bram_07_INIT_12,
    INIT_13 => rom_bram_07_INIT_13,
    INIT_14 => rom_bram_07_INIT_14,
    INIT_15 => rom_bram_07_INIT_15,
    INIT_16 => rom_bram_07_INIT_16,
    INIT_17 => rom_bram_07_INIT_17,
    INIT_18 => rom_bram_07_INIT_18,
    INIT_19 => rom_bram_07_INIT_19,
    INIT_1A => rom_bram_07_INIT_1A,
    INIT_1B => rom_bram_07_INIT_1B,
    INIT_1C => rom_bram_07_INIT_1C,
    INIT_1D => rom_bram_07_INIT_1D,
    INIT_1E => rom_bram_07_INIT_1E,
    INIT_1F => rom_bram_07_INIT_1F,
    INIT_20 => rom_bram_07_INIT_20,
    INIT_21 => rom_bram_07_INIT_21,
    INIT_22 => rom_bram_07_INIT_22,
    INIT_23 => rom_bram_07_INIT_23,
    INIT_24 => rom_bram_07_INIT_24,
    INIT_25 => rom_bram_07_INIT_25,
    INIT_26 => rom_bram_07_INIT_26,
    INIT_27 => rom_bram_07_INIT_27,
    INIT_28 => rom_bram_07_INIT_28,
    INIT_29 => rom_bram_07_INIT_29,
    INIT_2A => rom_bram_07_INIT_2A,
    INIT_2B => rom_bram_07_INIT_2B,
    INIT_2C => rom_bram_07_INIT_2C,
    INIT_2D => rom_bram_07_INIT_2D,
    INIT_2E => rom_bram_07_INIT_2E,
    INIT_2F => rom_bram_07_INIT_2F,
    INIT_30 => rom_bram_07_INIT_30,
    INIT_31 => rom_bram_07_INIT_31,
    INIT_32 => rom_bram_07_INIT_32,
    INIT_33 => rom_bram_07_INIT_33,
    INIT_34 => rom_bram_07_INIT_34,
    INIT_35 => rom_bram_07_INIT_35,
    INIT_36 => rom_bram_07_INIT_36,
    INIT_37 => rom_bram_07_INIT_37,
    INIT_38 => rom_bram_07_INIT_38,
    INIT_39 => rom_bram_07_INIT_39,
    INIT_3A => rom_bram_07_INIT_3A,
    INIT_3B => rom_bram_07_INIT_3B,
    INIT_3C => rom_bram_07_INIT_3C,
    INIT_3D => rom_bram_07_INIT_3D,
    INIT_3E => rom_bram_07_INIT_3E,
    INIT_3F => rom_bram_07_INIT_3F )
  PORT MAP( 
    DO => rom_bram_07_dat_o,
    dop => OPEN,    
    di => "00000000",
    dip => "0",
    addr => adr_i(10 DOWNTO 0), 
    clk => clk_i,    
    en => '1',
    ssr => '0',
    we => '0' );

  -- BRAM 8 in address space [0x00004000:0x000047FF], bit lane [7:0]
  rom_bram_08 : RAMB16_S9 
  GENERIC MAP(
    INIT_00 => rom_bram_08_INIT_00,
    INIT_01 => rom_bram_08_INIT_01,
    INIT_02 => rom_bram_08_INIT_02,
    INIT_03 => rom_bram_08_INIT_03,
    INIT_04 => rom_bram_08_INIT_04,
    INIT_05 => rom_bram_08_INIT_05,
    INIT_06 => rom_bram_08_INIT_06,
    INIT_07 => rom_bram_08_INIT_07,
    INIT_08 => rom_bram_08_INIT_08,
    INIT_09 => rom_bram_08_INIT_09,
    INIT_0A => rom_bram_08_INIT_0A,
    INIT_0B => rom_bram_08_INIT_0B,
    INIT_0C => rom_bram_08_INIT_0C,
    INIT_0D => rom_bram_08_INIT_0D,
    INIT_0E => rom_bram_08_INIT_0E,
    INIT_0F => rom_bram_08_INIT_0F,
    INIT_10 => rom_bram_08_INIT_10,
    INIT_11 => rom_bram_08_INIT_11,
    INIT_12 => rom_bram_08_INIT_12,
    INIT_13 => rom_bram_08_INIT_13,
    INIT_14 => rom_bram_08_INIT_14,
    INIT_15 => rom_bram_08_INIT_15,
    INIT_16 => rom_bram_08_INIT_16,
    INIT_17 => rom_bram_08_INIT_17,
    INIT_18 => rom_bram_08_INIT_18,
    INIT_19 => rom_bram_08_INIT_19,
    INIT_1A => rom_bram_08_INIT_1A,
    INIT_1B => rom_bram_08_INIT_1B,
    INIT_1C => rom_bram_08_INIT_1C,
    INIT_1D => rom_bram_08_INIT_1D,
    INIT_1E => rom_bram_08_INIT_1E,
    INIT_1F => rom_bram_08_INIT_1F,
    INIT_20 => rom_bram_08_INIT_20,
    INIT_21 => rom_bram_08_INIT_21,
    INIT_22 => rom_bram_08_INIT_22,
    INIT_23 => rom_bram_08_INIT_23,
    INIT_24 => rom_bram_08_INIT_24,
    INIT_25 => rom_bram_08_INIT_25,
    INIT_26 => rom_bram_08_INIT_26,
    INIT_27 => rom_bram_08_INIT_27,
    INIT_28 => rom_bram_08_INIT_28,
    INIT_29 => rom_bram_08_INIT_29,
    INIT_2A => rom_bram_08_INIT_2A,
    INIT_2B => rom_bram_08_INIT_2B,
    INIT_2C => rom_bram_08_INIT_2C,
    INIT_2D => rom_bram_08_INIT_2D,
    INIT_2E => rom_bram_08_INIT_2E,
    INIT_2F => rom_bram_08_INIT_2F,
    INIT_30 => rom_bram_08_INIT_30,
    INIT_31 => rom_bram_08_INIT_31,
    INIT_32 => rom_bram_08_INIT_32,
    INIT_33 => rom_bram_08_INIT_33,
    INIT_34 => rom_bram_08_INIT_34,
    INIT_35 => rom_bram_08_INIT_35,
    INIT_36 => rom_bram_08_INIT_36,
    INIT_37 => rom_bram_08_INIT_37,
    INIT_38 => rom_bram_08_INIT_38,
    INIT_39 => rom_bram_08_INIT_39,
    INIT_3A => rom_bram_08_INIT_3A,
    INIT_3B => rom_bram_08_INIT_3B,
    INIT_3C => rom_bram_08_INIT_3C,
    INIT_3D => rom_bram_08_INIT_3D,
    INIT_3E => rom_bram_08_INIT_3E,
    INIT_3F => rom_bram_08_INIT_3F )
  PORT MAP( 
    DO => rom_bram_08_dat_o,
    dop => OPEN,    
    di => "00000000",
    dip => "0",
    addr => adr_i(10 DOWNTO 0), 
    clk => clk_i,    
    en => '1',
    ssr => '0',
    we => '0' );

  -- BRAM 9 in address space [0x00004800:0x00004FFF], bit lane [7:0]
  rom_bram_09 : RAMB16_S9 
  GENERIC MAP(
    INIT_00 => rom_bram_09_INIT_00,
    INIT_01 => rom_bram_09_INIT_01,
    INIT_02 => rom_bram_09_INIT_02,
    INIT_03 => rom_bram_09_INIT_03,
    INIT_04 => rom_bram_09_INIT_04,
    INIT_05 => rom_bram_09_INIT_05,
    INIT_06 => rom_bram_09_INIT_06,
    INIT_07 => rom_bram_09_INIT_07,
    INIT_08 => rom_bram_09_INIT_08,
    INIT_09 => rom_bram_09_INIT_09,
    INIT_0A => rom_bram_09_INIT_0A,
    INIT_0B => rom_bram_09_INIT_0B,
    INIT_0C => rom_bram_09_INIT_0C,
    INIT_0D => rom_bram_09_INIT_0D,
    INIT_0E => rom_bram_09_INIT_0E,
    INIT_0F => rom_bram_09_INIT_0F,
    INIT_10 => rom_bram_09_INIT_10,
    INIT_11 => rom_bram_09_INIT_11,
    INIT_12 => rom_bram_09_INIT_12,
    INIT_13 => rom_bram_09_INIT_13,
    INIT_14 => rom_bram_09_INIT_14,
    INIT_15 => rom_bram_09_INIT_15,
    INIT_16 => rom_bram_09_INIT_16,
    INIT_17 => rom_bram_09_INIT_17,
    INIT_18 => rom_bram_09_INIT_18,
    INIT_19 => rom_bram_09_INIT_19,
    INIT_1A => rom_bram_09_INIT_1A,
    INIT_1B => rom_bram_09_INIT_1B,
    INIT_1C => rom_bram_09_INIT_1C,
    INIT_1D => rom_bram_09_INIT_1D,
    INIT_1E => rom_bram_09_INIT_1E,
    INIT_1F => rom_bram_09_INIT_1F,
    INIT_20 => rom_bram_09_INIT_20,
    INIT_21 => rom_bram_09_INIT_21,
    INIT_22 => rom_bram_09_INIT_22,
    INIT_23 => rom_bram_09_INIT_23,
    INIT_24 => rom_bram_09_INIT_24,
    INIT_25 => rom_bram_09_INIT_25,
    INIT_26 => rom_bram_09_INIT_26,
    INIT_27 => rom_bram_09_INIT_27,
    INIT_28 => rom_bram_09_INIT_28,
    INIT_29 => rom_bram_09_INIT_29,
    INIT_2A => rom_bram_09_INIT_2A,
    INIT_2B => rom_bram_09_INIT_2B,
    INIT_2C => rom_bram_09_INIT_2C,
    INIT_2D => rom_bram_09_INIT_2D,
    INIT_2E => rom_bram_09_INIT_2E,
    INIT_2F => rom_bram_09_INIT_2F,
    INIT_30 => rom_bram_09_INIT_30,
    INIT_31 => rom_bram_09_INIT_31,
    INIT_32 => rom_bram_09_INIT_32,
    INIT_33 => rom_bram_09_INIT_33,
    INIT_34 => rom_bram_09_INIT_34,
    INIT_35 => rom_bram_09_INIT_35,
    INIT_36 => rom_bram_09_INIT_36,
    INIT_37 => rom_bram_09_INIT_37,
    INIT_38 => rom_bram_09_INIT_38,
    INIT_39 => rom_bram_09_INIT_39,
    INIT_3A => rom_bram_09_INIT_3A,
    INIT_3B => rom_bram_09_INIT_3B,
    INIT_3C => rom_bram_09_INIT_3C,
    INIT_3D => rom_bram_09_INIT_3D,
    INIT_3E => rom_bram_09_INIT_3E,
    INIT_3F => rom_bram_09_INIT_3F )
  PORT MAP( 
    DO => rom_bram_09_dat_o,
    dop => OPEN,    
    di => "00000000",
    dip => "0",
    addr => adr_i(10 DOWNTO 0), 
    clk => clk_i,    
    en => '1',
    ssr => '0',
    we => '0' );
    
  -- BRAM A in address space [0x00005000:0x000057FF], bit lane [7:0]
  rom_bram_0A : RAMB16_S9 
  GENERIC MAP(
    INIT_00 => rom_bram_0A_INIT_00,
    INIT_01 => rom_bram_0A_INIT_01,
    INIT_02 => rom_bram_0A_INIT_02,
    INIT_03 => rom_bram_0A_INIT_03,
    INIT_04 => rom_bram_0A_INIT_04,
    INIT_05 => rom_bram_0A_INIT_05,
    INIT_06 => rom_bram_0A_INIT_06,
    INIT_07 => rom_bram_0A_INIT_07,
    INIT_08 => rom_bram_0A_INIT_08,
    INIT_09 => rom_bram_0A_INIT_09,
    INIT_0A => rom_bram_0A_INIT_0A,
    INIT_0B => rom_bram_0A_INIT_0B,
    INIT_0C => rom_bram_0A_INIT_0C,
    INIT_0D => rom_bram_0A_INIT_0D,
    INIT_0E => rom_bram_0A_INIT_0E,
    INIT_0F => rom_bram_0A_INIT_0F,
    INIT_10 => rom_bram_0A_INIT_10,
    INIT_11 => rom_bram_0A_INIT_11,
    INIT_12 => rom_bram_0A_INIT_12,
    INIT_13 => rom_bram_0A_INIT_13,
    INIT_14 => rom_bram_0A_INIT_14,
    INIT_15 => rom_bram_0A_INIT_15,
    INIT_16 => rom_bram_0A_INIT_16,
    INIT_17 => rom_bram_0A_INIT_17,
    INIT_18 => rom_bram_0A_INIT_18,
    INIT_19 => rom_bram_0A_INIT_19,
    INIT_1A => rom_bram_0A_INIT_1A,
    INIT_1B => rom_bram_0A_INIT_1B,
    INIT_1C => rom_bram_0A_INIT_1C,
    INIT_1D => rom_bram_0A_INIT_1D,
    INIT_1E => rom_bram_0A_INIT_1E,
    INIT_1F => rom_bram_0A_INIT_1F,
    INIT_20 => rom_bram_0A_INIT_20,
    INIT_21 => rom_bram_0A_INIT_21,
    INIT_22 => rom_bram_0A_INIT_22,
    INIT_23 => rom_bram_0A_INIT_23,
    INIT_24 => rom_bram_0A_INIT_24,
    INIT_25 => rom_bram_0A_INIT_25,
    INIT_26 => rom_bram_0A_INIT_26,
    INIT_27 => rom_bram_0A_INIT_27,
    INIT_28 => rom_bram_0A_INIT_28,
    INIT_29 => rom_bram_0A_INIT_29,
    INIT_2A => rom_bram_0A_INIT_2A,
    INIT_2B => rom_bram_0A_INIT_2B,
    INIT_2C => rom_bram_0A_INIT_2C,
    INIT_2D => rom_bram_0A_INIT_2D,
    INIT_2E => rom_bram_0A_INIT_2E,
    INIT_2F => rom_bram_0A_INIT_2F,
    INIT_30 => rom_bram_0A_INIT_30,
    INIT_31 => rom_bram_0A_INIT_31,
    INIT_32 => rom_bram_0A_INIT_32,
    INIT_33 => rom_bram_0A_INIT_33,
    INIT_34 => rom_bram_0A_INIT_34,
    INIT_35 => rom_bram_0A_INIT_35,
    INIT_36 => rom_bram_0A_INIT_36,
    INIT_37 => rom_bram_0A_INIT_37,
    INIT_38 => rom_bram_0A_INIT_38,
    INIT_39 => rom_bram_0A_INIT_39,
    INIT_3A => rom_bram_0A_INIT_3A,
    INIT_3B => rom_bram_0A_INIT_3B,
    INIT_3C => rom_bram_0A_INIT_3C,
    INIT_3D => rom_bram_0A_INIT_3D,
    INIT_3E => rom_bram_0A_INIT_3E,
    INIT_3F => rom_bram_0A_INIT_3F )
  PORT MAP( 
    DO => rom_bram_0A_dat_o,
    dop => OPEN,    
    di => "00000000",
    dip => "0",
    addr => adr_i(10 DOWNTO 0), 
    clk => clk_i,    
    en => '1',
    ssr => '0',
    we => '0' );
    
  -- BRAM B in address space [0x00005800:0x00005FFF], bit lane [7:0]
  rom_bram_0B : RAMB16_S9 
  GENERIC MAP(
    INIT_00 => rom_bram_0B_INIT_00,
    INIT_01 => rom_bram_0B_INIT_01,
    INIT_02 => rom_bram_0B_INIT_02,
    INIT_03 => rom_bram_0B_INIT_03,
    INIT_04 => rom_bram_0B_INIT_04,
    INIT_05 => rom_bram_0B_INIT_05,
    INIT_06 => rom_bram_0B_INIT_06,
    INIT_07 => rom_bram_0B_INIT_07,
    INIT_08 => rom_bram_0B_INIT_08,
    INIT_09 => rom_bram_0B_INIT_09,
    INIT_0A => rom_bram_0B_INIT_0A,
    INIT_0B => rom_bram_0B_INIT_0B,
    INIT_0C => rom_bram_0B_INIT_0C,
    INIT_0D => rom_bram_0B_INIT_0D,
    INIT_0E => rom_bram_0B_INIT_0E,
    INIT_0F => rom_bram_0B_INIT_0F,
    INIT_10 => rom_bram_0B_INIT_10,
    INIT_11 => rom_bram_0B_INIT_11,
    INIT_12 => rom_bram_0B_INIT_12,
    INIT_13 => rom_bram_0B_INIT_13,
    INIT_14 => rom_bram_0B_INIT_14,
    INIT_15 => rom_bram_0B_INIT_15,
    INIT_16 => rom_bram_0B_INIT_16,
    INIT_17 => rom_bram_0B_INIT_17,
    INIT_18 => rom_bram_0B_INIT_18,
    INIT_19 => rom_bram_0B_INIT_19,
    INIT_1A => rom_bram_0B_INIT_1A,
    INIT_1B => rom_bram_0B_INIT_1B,
    INIT_1C => rom_bram_0B_INIT_1C,
    INIT_1D => rom_bram_0B_INIT_1D,
    INIT_1E => rom_bram_0B_INIT_1E,
    INIT_1F => rom_bram_0B_INIT_1F,
    INIT_20 => rom_bram_0B_INIT_20,
    INIT_21 => rom_bram_0B_INIT_21,
    INIT_22 => rom_bram_0B_INIT_22,
    INIT_23 => rom_bram_0B_INIT_23,
    INIT_24 => rom_bram_0B_INIT_24,
    INIT_25 => rom_bram_0B_INIT_25,
    INIT_26 => rom_bram_0B_INIT_26,
    INIT_27 => rom_bram_0B_INIT_27,
    INIT_28 => rom_bram_0B_INIT_28,
    INIT_29 => rom_bram_0B_INIT_29,
    INIT_2A => rom_bram_0B_INIT_2A,
    INIT_2B => rom_bram_0B_INIT_2B,
    INIT_2C => rom_bram_0B_INIT_2C,
    INIT_2D => rom_bram_0B_INIT_2D,
    INIT_2E => rom_bram_0B_INIT_2E,
    INIT_2F => rom_bram_0B_INIT_2F,
    INIT_30 => rom_bram_0B_INIT_30,
    INIT_31 => rom_bram_0B_INIT_31,
    INIT_32 => rom_bram_0B_INIT_32,
    INIT_33 => rom_bram_0B_INIT_33,
    INIT_34 => rom_bram_0B_INIT_34,
    INIT_35 => rom_bram_0B_INIT_35,
    INIT_36 => rom_bram_0B_INIT_36,
    INIT_37 => rom_bram_0B_INIT_37,
    INIT_38 => rom_bram_0B_INIT_38,
    INIT_39 => rom_bram_0B_INIT_39,
    INIT_3A => rom_bram_0B_INIT_3A,
    INIT_3B => rom_bram_0B_INIT_3B,
    INIT_3C => rom_bram_0B_INIT_3C,
    INIT_3D => rom_bram_0B_INIT_3D,
    INIT_3E => rom_bram_0B_INIT_3E,
    INIT_3F => rom_bram_0B_INIT_3F )
  PORT MAP( 
    DO => rom_bram_0B_dat_o,
    dop => OPEN,    
    di => "00000000",
    dip => "0",
    addr => adr_i(10 DOWNTO 0), 
    clk => clk_i,    
    en => '1',
    ssr => '0',
    we => '0' ); 
  
  -- BRAM C in address space [0x00006000:0x000067FF], bit lane [7:0]
  rom_bram_0C : RAMB16_S9 
  GENERIC MAP(
    INIT_00 => rom_bram_0C_INIT_00,
    INIT_01 => rom_bram_0C_INIT_01,
    INIT_02 => rom_bram_0C_INIT_02,
    INIT_03 => rom_bram_0C_INIT_03,
    INIT_04 => rom_bram_0C_INIT_04,
    INIT_05 => rom_bram_0C_INIT_05,
    INIT_06 => rom_bram_0C_INIT_06,
    INIT_07 => rom_bram_0C_INIT_07,
    INIT_08 => rom_bram_0C_INIT_08,
    INIT_09 => rom_bram_0C_INIT_09,
    INIT_0A => rom_bram_0C_INIT_0A,
    INIT_0B => rom_bram_0C_INIT_0B,
    INIT_0C => rom_bram_0C_INIT_0C,
    INIT_0D => rom_bram_0C_INIT_0D,
    INIT_0E => rom_bram_0C_INIT_0E,
    INIT_0F => rom_bram_0C_INIT_0F,
    INIT_10 => rom_bram_0C_INIT_10,
    INIT_11 => rom_bram_0C_INIT_11,
    INIT_12 => rom_bram_0C_INIT_12,
    INIT_13 => rom_bram_0C_INIT_13,
    INIT_14 => rom_bram_0C_INIT_14,
    INIT_15 => rom_bram_0C_INIT_15,
    INIT_16 => rom_bram_0C_INIT_16,
    INIT_17 => rom_bram_0C_INIT_17,
    INIT_18 => rom_bram_0C_INIT_18,
    INIT_19 => rom_bram_0C_INIT_19,
    INIT_1A => rom_bram_0C_INIT_1A,
    INIT_1B => rom_bram_0C_INIT_1B,
    INIT_1C => rom_bram_0C_INIT_1C,
    INIT_1D => rom_bram_0C_INIT_1D,
    INIT_1E => rom_bram_0C_INIT_1E,
    INIT_1F => rom_bram_0C_INIT_1F,
    INIT_20 => rom_bram_0C_INIT_20,
    INIT_21 => rom_bram_0C_INIT_21,
    INIT_22 => rom_bram_0C_INIT_22,
    INIT_23 => rom_bram_0C_INIT_23,
    INIT_24 => rom_bram_0C_INIT_24,
    INIT_25 => rom_bram_0C_INIT_25,
    INIT_26 => rom_bram_0C_INIT_26,
    INIT_27 => rom_bram_0C_INIT_27,
    INIT_28 => rom_bram_0C_INIT_28,
    INIT_29 => rom_bram_0C_INIT_29,
    INIT_2A => rom_bram_0C_INIT_2A,
    INIT_2B => rom_bram_0C_INIT_2B,
    INIT_2C => rom_bram_0C_INIT_2C,
    INIT_2D => rom_bram_0C_INIT_2D,
    INIT_2E => rom_bram_0C_INIT_2E,
    INIT_2F => rom_bram_0C_INIT_2F,
    INIT_30 => rom_bram_0C_INIT_30,
    INIT_31 => rom_bram_0C_INIT_31,
    INIT_32 => rom_bram_0C_INIT_32,
    INIT_33 => rom_bram_0C_INIT_33,
    INIT_34 => rom_bram_0C_INIT_34,
    INIT_35 => rom_bram_0C_INIT_35,
    INIT_36 => rom_bram_0C_INIT_36,
    INIT_37 => rom_bram_0C_INIT_37,
    INIT_38 => rom_bram_0C_INIT_38,
    INIT_39 => rom_bram_0C_INIT_39,
    INIT_3A => rom_bram_0C_INIT_3A,
    INIT_3B => rom_bram_0C_INIT_3B,
    INIT_3C => rom_bram_0C_INIT_3C,
    INIT_3D => rom_bram_0C_INIT_3D,
    INIT_3E => rom_bram_0C_INIT_3E,
    INIT_3F => rom_bram_0C_INIT_3F )
  PORT MAP( 
    DO => rom_bram_0C_dat_o,
    dop => OPEN,    
    di => "00000000",
    dip => "0",
    addr => adr_i(10 DOWNTO 0), 
    clk => clk_i,    
    en => '1',
    ssr => '0',
    we => '0' );

  -- BRAM D in address space [0x00006800:0x00006FFF], bit lane [7:0]
  rom_bram_0D : RAMB16_S9 
  GENERIC MAP(
    INIT_00 => rom_bram_0D_INIT_00,
    INIT_01 => rom_bram_0D_INIT_01,
    INIT_02 => rom_bram_0D_INIT_02,
    INIT_03 => rom_bram_0D_INIT_03,
    INIT_04 => rom_bram_0D_INIT_04,
    INIT_05 => rom_bram_0D_INIT_05,
    INIT_06 => rom_bram_0D_INIT_06,
    INIT_07 => rom_bram_0D_INIT_07,
    INIT_08 => rom_bram_0D_INIT_08,
    INIT_09 => rom_bram_0D_INIT_09,
    INIT_0A => rom_bram_0D_INIT_0A,
    INIT_0B => rom_bram_0D_INIT_0B,
    INIT_0C => rom_bram_0D_INIT_0C,
    INIT_0D => rom_bram_0D_INIT_0D,
    INIT_0E => rom_bram_0D_INIT_0E,
    INIT_0F => rom_bram_0D_INIT_0F,
    INIT_10 => rom_bram_0D_INIT_10,
    INIT_11 => rom_bram_0D_INIT_11,
    INIT_12 => rom_bram_0D_INIT_12,
    INIT_13 => rom_bram_0D_INIT_13,
    INIT_14 => rom_bram_0D_INIT_14,
    INIT_15 => rom_bram_0D_INIT_15,
    INIT_16 => rom_bram_0D_INIT_16,
    INIT_17 => rom_bram_0D_INIT_17,
    INIT_18 => rom_bram_0D_INIT_18,
    INIT_19 => rom_bram_0D_INIT_19,
    INIT_1A => rom_bram_0D_INIT_1A,
    INIT_1B => rom_bram_0D_INIT_1B,
    INIT_1C => rom_bram_0D_INIT_1C,
    INIT_1D => rom_bram_0D_INIT_1D,
    INIT_1E => rom_bram_0D_INIT_1E,
    INIT_1F => rom_bram_0D_INIT_1F,
    INIT_20 => rom_bram_0D_INIT_20,
    INIT_21 => rom_bram_0D_INIT_21,
    INIT_22 => rom_bram_0D_INIT_22,
    INIT_23 => rom_bram_0D_INIT_23,
    INIT_24 => rom_bram_0D_INIT_24,
    INIT_25 => rom_bram_0D_INIT_25,
    INIT_26 => rom_bram_0D_INIT_26,
    INIT_27 => rom_bram_0D_INIT_27,
    INIT_28 => rom_bram_0D_INIT_28,
    INIT_29 => rom_bram_0D_INIT_29,
    INIT_2A => rom_bram_0D_INIT_2A,
    INIT_2B => rom_bram_0D_INIT_2B,
    INIT_2C => rom_bram_0D_INIT_2C,
    INIT_2D => rom_bram_0D_INIT_2D,
    INIT_2E => rom_bram_0D_INIT_2E,
    INIT_2F => rom_bram_0D_INIT_2F,
    INIT_30 => rom_bram_0D_INIT_30,
    INIT_31 => rom_bram_0D_INIT_31,
    INIT_32 => rom_bram_0D_INIT_32,
    INIT_33 => rom_bram_0D_INIT_33,
    INIT_34 => rom_bram_0D_INIT_34,
    INIT_35 => rom_bram_0D_INIT_35,
    INIT_36 => rom_bram_0D_INIT_36,
    INIT_37 => rom_bram_0D_INIT_37,
    INIT_38 => rom_bram_0D_INIT_38,
    INIT_39 => rom_bram_0D_INIT_39,
    INIT_3A => rom_bram_0D_INIT_3A,
    INIT_3B => rom_bram_0D_INIT_3B,
    INIT_3C => rom_bram_0D_INIT_3C,
    INIT_3D => rom_bram_0D_INIT_3D,
    INIT_3E => rom_bram_0D_INIT_3E,
    INIT_3F => rom_bram_0D_INIT_3F )
  PORT MAP( 
    DO => rom_bram_0D_dat_o,
    dop => OPEN,    
    di => "00000000",
    dip => "0",
    addr => adr_i(10 DOWNTO 0), 
    clk => clk_i,    
    en => '1',
    ssr => '0',
    we => '0' );
    
  -- BRAM E in address space [0x00007000:0x000077FF], bit lane [7:0]
  rom_bram_0E : RAMB16_S9 
  GENERIC MAP(
    INIT_00 => rom_bram_0E_INIT_00,
    INIT_01 => rom_bram_0E_INIT_01,
    INIT_02 => rom_bram_0E_INIT_02,
    INIT_03 => rom_bram_0E_INIT_03,
    INIT_04 => rom_bram_0E_INIT_04,
    INIT_05 => rom_bram_0E_INIT_05,
    INIT_06 => rom_bram_0E_INIT_06,
    INIT_07 => rom_bram_0E_INIT_07,
    INIT_08 => rom_bram_0E_INIT_08,
    INIT_09 => rom_bram_0E_INIT_09,
    INIT_0A => rom_bram_0E_INIT_0A,
    INIT_0B => rom_bram_0E_INIT_0B,
    INIT_0C => rom_bram_0E_INIT_0C,
    INIT_0D => rom_bram_0E_INIT_0D,
    INIT_0E => rom_bram_0E_INIT_0E,
    INIT_0F => rom_bram_0E_INIT_0F,
    INIT_10 => rom_bram_0E_INIT_10,
    INIT_11 => rom_bram_0E_INIT_11,
    INIT_12 => rom_bram_0E_INIT_12,
    INIT_13 => rom_bram_0E_INIT_13,
    INIT_14 => rom_bram_0E_INIT_14,
    INIT_15 => rom_bram_0E_INIT_15,
    INIT_16 => rom_bram_0E_INIT_16,
    INIT_17 => rom_bram_0E_INIT_17,
    INIT_18 => rom_bram_0E_INIT_18,
    INIT_19 => rom_bram_0E_INIT_19,
    INIT_1A => rom_bram_0E_INIT_1A,
    INIT_1B => rom_bram_0E_INIT_1B,
    INIT_1C => rom_bram_0E_INIT_1C,
    INIT_1D => rom_bram_0E_INIT_1D,
    INIT_1E => rom_bram_0E_INIT_1E,
    INIT_1F => rom_bram_0E_INIT_1F,
    INIT_20 => rom_bram_0E_INIT_20,
    INIT_21 => rom_bram_0E_INIT_21,
    INIT_22 => rom_bram_0E_INIT_22,
    INIT_23 => rom_bram_0E_INIT_23,
    INIT_24 => rom_bram_0E_INIT_24,
    INIT_25 => rom_bram_0E_INIT_25,
    INIT_26 => rom_bram_0E_INIT_26,
    INIT_27 => rom_bram_0E_INIT_27,
    INIT_28 => rom_bram_0E_INIT_28,
    INIT_29 => rom_bram_0E_INIT_29,
    INIT_2A => rom_bram_0E_INIT_2A,
    INIT_2B => rom_bram_0E_INIT_2B,
    INIT_2C => rom_bram_0E_INIT_2C,
    INIT_2D => rom_bram_0E_INIT_2D,
    INIT_2E => rom_bram_0E_INIT_2E,
    INIT_2F => rom_bram_0E_INIT_2F,
    INIT_30 => rom_bram_0E_INIT_30,
    INIT_31 => rom_bram_0E_INIT_31,
    INIT_32 => rom_bram_0E_INIT_32,
    INIT_33 => rom_bram_0E_INIT_33,
    INIT_34 => rom_bram_0E_INIT_34,
    INIT_35 => rom_bram_0E_INIT_35,
    INIT_36 => rom_bram_0E_INIT_36,
    INIT_37 => rom_bram_0E_INIT_37,
    INIT_38 => rom_bram_0E_INIT_38,
    INIT_39 => rom_bram_0E_INIT_39,
    INIT_3A => rom_bram_0E_INIT_3A,
    INIT_3B => rom_bram_0E_INIT_3B,
    INIT_3C => rom_bram_0E_INIT_3C,
    INIT_3D => rom_bram_0E_INIT_3D,
    INIT_3E => rom_bram_0E_INIT_3E,
    INIT_3F => rom_bram_0E_INIT_3F )
  PORT MAP( 
    DO => rom_bram_0E_dat_o,
    dop => OPEN,    
    di => "00000000",
    dip => "0",
    addr => adr_i(10 DOWNTO 0), 
    clk => clk_i,    
    en => '1',
    ssr => '0',
    we => '0' );
    
  -- BRAM F in address space [0x00007800:0x00007FFF], bit lane [7:0]
  rom_bram_0F : RAMB16_S9 
  GENERIC MAP(
    INIT_00 => rom_bram_0F_INIT_00,
    INIT_01 => rom_bram_0F_INIT_01,
    INIT_02 => rom_bram_0F_INIT_02,
    INIT_03 => rom_bram_0F_INIT_03,
    INIT_04 => rom_bram_0F_INIT_04,
    INIT_05 => rom_bram_0F_INIT_05,
    INIT_06 => rom_bram_0F_INIT_06,
    INIT_07 => rom_bram_0F_INIT_07,
    INIT_08 => rom_bram_0F_INIT_08,
    INIT_09 => rom_bram_0F_INIT_09,
    INIT_0A => rom_bram_0F_INIT_0A,
    INIT_0B => rom_bram_0F_INIT_0B,
    INIT_0C => rom_bram_0F_INIT_0C,
    INIT_0D => rom_bram_0F_INIT_0D,
    INIT_0E => rom_bram_0F_INIT_0E,
    INIT_0F => rom_bram_0F_INIT_0F,
    INIT_10 => rom_bram_0F_INIT_10,
    INIT_11 => rom_bram_0F_INIT_11,
    INIT_12 => rom_bram_0F_INIT_12,
    INIT_13 => rom_bram_0F_INIT_13,
    INIT_14 => rom_bram_0F_INIT_14,
    INIT_15 => rom_bram_0F_INIT_15,
    INIT_16 => rom_bram_0F_INIT_16,
    INIT_17 => rom_bram_0F_INIT_17,
    INIT_18 => rom_bram_0F_INIT_18,
    INIT_19 => rom_bram_0F_INIT_19,
    INIT_1A => rom_bram_0F_INIT_1A,
    INIT_1B => rom_bram_0F_INIT_1B,
    INIT_1C => rom_bram_0F_INIT_1C,
    INIT_1D => rom_bram_0F_INIT_1D,
    INIT_1E => rom_bram_0F_INIT_1E,
    INIT_1F => rom_bram_0F_INIT_1F,
    INIT_20 => rom_bram_0F_INIT_20,
    INIT_21 => rom_bram_0F_INIT_21,
    INIT_22 => rom_bram_0F_INIT_22,
    INIT_23 => rom_bram_0F_INIT_23,
    INIT_24 => rom_bram_0F_INIT_24,
    INIT_25 => rom_bram_0F_INIT_25,
    INIT_26 => rom_bram_0F_INIT_26,
    INIT_27 => rom_bram_0F_INIT_27,
    INIT_28 => rom_bram_0F_INIT_28,
    INIT_29 => rom_bram_0F_INIT_29,
    INIT_2A => rom_bram_0F_INIT_2A,
    INIT_2B => rom_bram_0F_INIT_2B,
    INIT_2C => rom_bram_0F_INIT_2C,
    INIT_2D => rom_bram_0F_INIT_2D,
    INIT_2E => rom_bram_0F_INIT_2E,
    INIT_2F => rom_bram_0F_INIT_2F,
    INIT_30 => rom_bram_0F_INIT_30,
    INIT_31 => rom_bram_0F_INIT_31,
    INIT_32 => rom_bram_0F_INIT_32,
    INIT_33 => rom_bram_0F_INIT_33,
    INIT_34 => rom_bram_0F_INIT_34,
    INIT_35 => rom_bram_0F_INIT_35,
    INIT_36 => rom_bram_0F_INIT_36,
    INIT_37 => rom_bram_0F_INIT_37,
    INIT_38 => rom_bram_0F_INIT_38,
    INIT_39 => rom_bram_0F_INIT_39,
    INIT_3A => rom_bram_0F_INIT_3A,
    INIT_3B => rom_bram_0F_INIT_3B,
    INIT_3C => rom_bram_0F_INIT_3C,
    INIT_3D => rom_bram_0F_INIT_3D,
    INIT_3E => rom_bram_0F_INIT_3E,
    INIT_3F => rom_bram_0F_INIT_3F )
  PORT MAP( 
    DO => rom_bram_0F_dat_o,
    dop => OPEN,    
    di => "00000000",
    dip => "0",
    addr => adr_i(10 DOWNTO 0), 
    clk => clk_i,    
    en => '1',
    ssr => '0',
    we => '0' );

  -- BRAM 10 in address space [0x00008000:0x000087FF], bit lane [7:0]
  rom_bram_10 : RAMB16_S9 
  GENERIC MAP(
    INIT_00 => rom_bram_10_INIT_00,
    INIT_01 => rom_bram_10_INIT_01,
    INIT_02 => rom_bram_10_INIT_02,
    INIT_03 => rom_bram_10_INIT_03,
    INIT_04 => rom_bram_10_INIT_04,
    INIT_05 => rom_bram_10_INIT_05,
    INIT_06 => rom_bram_10_INIT_06,
    INIT_07 => rom_bram_10_INIT_07,
    INIT_08 => rom_bram_10_INIT_08,
    INIT_09 => rom_bram_10_INIT_09,
    INIT_0A => rom_bram_10_INIT_0A,
    INIT_0B => rom_bram_10_INIT_0B,
    INIT_0C => rom_bram_10_INIT_0C,
    INIT_0D => rom_bram_10_INIT_0D,
    INIT_0E => rom_bram_10_INIT_0E,
    INIT_0F => rom_bram_10_INIT_0F,
    INIT_10 => rom_bram_10_INIT_10,
    INIT_11 => rom_bram_10_INIT_11,
    INIT_12 => rom_bram_10_INIT_12,
    INIT_13 => rom_bram_10_INIT_13,
    INIT_14 => rom_bram_10_INIT_14,
    INIT_15 => rom_bram_10_INIT_15,
    INIT_16 => rom_bram_10_INIT_16,
    INIT_17 => rom_bram_10_INIT_17,
    INIT_18 => rom_bram_10_INIT_18,
    INIT_19 => rom_bram_10_INIT_19,
    INIT_1A => rom_bram_10_INIT_1A,
    INIT_1B => rom_bram_10_INIT_1B,
    INIT_1C => rom_bram_10_INIT_1C,
    INIT_1D => rom_bram_10_INIT_1D,
    INIT_1E => rom_bram_10_INIT_1E,
    INIT_1F => rom_bram_10_INIT_1F,
    INIT_20 => rom_bram_10_INIT_20,
    INIT_21 => rom_bram_10_INIT_21,
    INIT_22 => rom_bram_10_INIT_22,
    INIT_23 => rom_bram_10_INIT_23,
    INIT_24 => rom_bram_10_INIT_24,
    INIT_25 => rom_bram_10_INIT_25,
    INIT_26 => rom_bram_10_INIT_26,
    INIT_27 => rom_bram_10_INIT_27,
    INIT_28 => rom_bram_10_INIT_28,
    INIT_29 => rom_bram_10_INIT_29,
    INIT_2A => rom_bram_10_INIT_2A,
    INIT_2B => rom_bram_10_INIT_2B,
    INIT_2C => rom_bram_10_INIT_2C,
    INIT_2D => rom_bram_10_INIT_2D,
    INIT_2E => rom_bram_10_INIT_2E,
    INIT_2F => rom_bram_10_INIT_2F,
    INIT_30 => rom_bram_10_INIT_30,
    INIT_31 => rom_bram_10_INIT_31,
    INIT_32 => rom_bram_10_INIT_32,
    INIT_33 => rom_bram_10_INIT_33,
    INIT_34 => rom_bram_10_INIT_34,
    INIT_35 => rom_bram_10_INIT_35,
    INIT_36 => rom_bram_10_INIT_36,
    INIT_37 => rom_bram_10_INIT_37,
    INIT_38 => rom_bram_10_INIT_38,
    INIT_39 => rom_bram_10_INIT_39,
    INIT_3A => rom_bram_10_INIT_3A,
    INIT_3B => rom_bram_10_INIT_3B,
    INIT_3C => rom_bram_10_INIT_3C,
    INIT_3D => rom_bram_10_INIT_3D,
    INIT_3E => rom_bram_10_INIT_3E,
    INIT_3F => rom_bram_10_INIT_3F )
  PORT MAP( 
    DO => rom_bram_10_dat_o,
    dop => OPEN,    
    di => "00000000",
    dip => "0",
    addr => adr_i(10 DOWNTO 0), 
    clk => clk_i,    
    en => '1',
    ssr => '0',
    we => '0' );

  -- BRAM 11 in address space [0x00008800:0x00008FFF], bit lane [7:0]
  rom_bram_11 : RAMB16_S9 
  GENERIC MAP(
    INIT_00 => rom_bram_11_INIT_00,
    INIT_01 => rom_bram_11_INIT_01,
    INIT_02 => rom_bram_11_INIT_02,
    INIT_03 => rom_bram_11_INIT_03,
    INIT_04 => rom_bram_11_INIT_04,
    INIT_05 => rom_bram_11_INIT_05,
    INIT_06 => rom_bram_11_INIT_06,
    INIT_07 => rom_bram_11_INIT_07,
    INIT_08 => rom_bram_11_INIT_08,
    INIT_09 => rom_bram_11_INIT_09,
    INIT_0A => rom_bram_11_INIT_0A,
    INIT_0B => rom_bram_11_INIT_0B,
    INIT_0C => rom_bram_11_INIT_0C,
    INIT_0D => rom_bram_11_INIT_0D,
    INIT_0E => rom_bram_11_INIT_0E,
    INIT_0F => rom_bram_11_INIT_0F,
    INIT_10 => rom_bram_11_INIT_10,
    INIT_11 => rom_bram_11_INIT_11,
    INIT_12 => rom_bram_11_INIT_12,
    INIT_13 => rom_bram_11_INIT_13,
    INIT_14 => rom_bram_11_INIT_14,
    INIT_15 => rom_bram_11_INIT_15,
    INIT_16 => rom_bram_11_INIT_16,
    INIT_17 => rom_bram_11_INIT_17,
    INIT_18 => rom_bram_11_INIT_18,
    INIT_19 => rom_bram_11_INIT_19,
    INIT_1A => rom_bram_11_INIT_1A,
    INIT_1B => rom_bram_11_INIT_1B,
    INIT_1C => rom_bram_11_INIT_1C,
    INIT_1D => rom_bram_11_INIT_1D,
    INIT_1E => rom_bram_11_INIT_1E,
    INIT_1F => rom_bram_11_INIT_1F,
    INIT_20 => rom_bram_11_INIT_20,
    INIT_21 => rom_bram_11_INIT_21,
    INIT_22 => rom_bram_11_INIT_22,
    INIT_23 => rom_bram_11_INIT_23,
    INIT_24 => rom_bram_11_INIT_24,
    INIT_25 => rom_bram_11_INIT_25,
    INIT_26 => rom_bram_11_INIT_26,
    INIT_27 => rom_bram_11_INIT_27,
    INIT_28 => rom_bram_11_INIT_28,
    INIT_29 => rom_bram_11_INIT_29,
    INIT_2A => rom_bram_11_INIT_2A,
    INIT_2B => rom_bram_11_INIT_2B,
    INIT_2C => rom_bram_11_INIT_2C,
    INIT_2D => rom_bram_11_INIT_2D,
    INIT_2E => rom_bram_11_INIT_2E,
    INIT_2F => rom_bram_11_INIT_2F,
    INIT_30 => rom_bram_11_INIT_30,
    INIT_31 => rom_bram_11_INIT_31,
    INIT_32 => rom_bram_11_INIT_32,
    INIT_33 => rom_bram_11_INIT_33,
    INIT_34 => rom_bram_11_INIT_34,
    INIT_35 => rom_bram_11_INIT_35,
    INIT_36 => rom_bram_11_INIT_36,
    INIT_37 => rom_bram_11_INIT_37,
    INIT_38 => rom_bram_11_INIT_38,
    INIT_39 => rom_bram_11_INIT_39,
    INIT_3A => rom_bram_11_INIT_3A,
    INIT_3B => rom_bram_11_INIT_3B,
    INIT_3C => rom_bram_11_INIT_3C,
    INIT_3D => rom_bram_11_INIT_3D,
    INIT_3E => rom_bram_11_INIT_3E,
    INIT_3F => rom_bram_11_INIT_3F )
  PORT MAP( 
    DO => rom_bram_11_dat_o,
    dop => OPEN,    
    di => "00000000",
    dip => "0",
    addr => adr_i(10 DOWNTO 0), 
    clk => clk_i,    
    en => '1',
    ssr => '0',
    we => '0' );
    
  -- BRAM 12 in address space [0x00009000:0x000097FF], bit lane [7:0]
  rom_bram_12 : RAMB16_S9 
  GENERIC MAP(
    INIT_00 => rom_bram_12_INIT_00,
    INIT_01 => rom_bram_12_INIT_01,
    INIT_02 => rom_bram_12_INIT_02,
    INIT_03 => rom_bram_12_INIT_03,
    INIT_04 => rom_bram_12_INIT_04,
    INIT_05 => rom_bram_12_INIT_05,
    INIT_06 => rom_bram_12_INIT_06,
    INIT_07 => rom_bram_12_INIT_07,
    INIT_08 => rom_bram_12_INIT_08,
    INIT_09 => rom_bram_12_INIT_09,
    INIT_0A => rom_bram_12_INIT_0A,
    INIT_0B => rom_bram_12_INIT_0B,
    INIT_0C => rom_bram_12_INIT_0C,
    INIT_0D => rom_bram_12_INIT_0D,
    INIT_0E => rom_bram_12_INIT_0E,
    INIT_0F => rom_bram_12_INIT_0F,
    INIT_10 => rom_bram_12_INIT_10,
    INIT_11 => rom_bram_12_INIT_11,
    INIT_12 => rom_bram_12_INIT_12,
    INIT_13 => rom_bram_12_INIT_13,
    INIT_14 => rom_bram_12_INIT_14,
    INIT_15 => rom_bram_12_INIT_15,
    INIT_16 => rom_bram_12_INIT_16,
    INIT_17 => rom_bram_12_INIT_17,
    INIT_18 => rom_bram_12_INIT_18,
    INIT_19 => rom_bram_12_INIT_19,
    INIT_1A => rom_bram_12_INIT_1A,
    INIT_1B => rom_bram_12_INIT_1B,
    INIT_1C => rom_bram_12_INIT_1C,
    INIT_1D => rom_bram_12_INIT_1D,
    INIT_1E => rom_bram_12_INIT_1E,
    INIT_1F => rom_bram_12_INIT_1F,
    INIT_20 => rom_bram_12_INIT_20,
    INIT_21 => rom_bram_12_INIT_21,
    INIT_22 => rom_bram_12_INIT_22,
    INIT_23 => rom_bram_12_INIT_23,
    INIT_24 => rom_bram_12_INIT_24,
    INIT_25 => rom_bram_12_INIT_25,
    INIT_26 => rom_bram_12_INIT_26,
    INIT_27 => rom_bram_12_INIT_27,
    INIT_28 => rom_bram_12_INIT_28,
    INIT_29 => rom_bram_12_INIT_29,
    INIT_2A => rom_bram_12_INIT_2A,
    INIT_2B => rom_bram_12_INIT_2B,
    INIT_2C => rom_bram_12_INIT_2C,
    INIT_2D => rom_bram_12_INIT_2D,
    INIT_2E => rom_bram_12_INIT_2E,
    INIT_2F => rom_bram_12_INIT_2F,
    INIT_30 => rom_bram_12_INIT_30,
    INIT_31 => rom_bram_12_INIT_31,
    INIT_32 => rom_bram_12_INIT_32,
    INIT_33 => rom_bram_12_INIT_33,
    INIT_34 => rom_bram_12_INIT_34,
    INIT_35 => rom_bram_12_INIT_35,
    INIT_36 => rom_bram_12_INIT_36,
    INIT_37 => rom_bram_12_INIT_37,
    INIT_38 => rom_bram_12_INIT_38,
    INIT_39 => rom_bram_12_INIT_39,
    INIT_3A => rom_bram_12_INIT_3A,
    INIT_3B => rom_bram_12_INIT_3B,
    INIT_3C => rom_bram_12_INIT_3C,
    INIT_3D => rom_bram_12_INIT_3D,
    INIT_3E => rom_bram_12_INIT_3E,
    INIT_3F => rom_bram_12_INIT_3F )
  PORT MAP( 
    DO => rom_bram_12_dat_o,
    dop => OPEN,    
    di => "00000000",
    dip => "0",
    addr => adr_i(10 DOWNTO 0), 
    clk => clk_i,    
    en => '1',
    ssr => '0',
    we => '0' );
    
  -- BRAM 13 in address space [0x00009800:0x00009FFF], bit lane [7:0]
  rom_bram_13 : RAMB16_S9 
  GENERIC MAP(
    INIT_00 => rom_bram_13_INIT_00,
    INIT_01 => rom_bram_13_INIT_01,
    INIT_02 => rom_bram_13_INIT_02,
    INIT_03 => rom_bram_13_INIT_03,
    INIT_04 => rom_bram_13_INIT_04,
    INIT_05 => rom_bram_13_INIT_05,
    INIT_06 => rom_bram_13_INIT_06,
    INIT_07 => rom_bram_13_INIT_07,
    INIT_08 => rom_bram_13_INIT_08,
    INIT_09 => rom_bram_13_INIT_09,
    INIT_0A => rom_bram_13_INIT_0A,
    INIT_0B => rom_bram_13_INIT_0B,
    INIT_0C => rom_bram_13_INIT_0C,
    INIT_0D => rom_bram_13_INIT_0D,
    INIT_0E => rom_bram_13_INIT_0E,
    INIT_0F => rom_bram_13_INIT_0F,
    INIT_10 => rom_bram_13_INIT_10,
    INIT_11 => rom_bram_13_INIT_11,
    INIT_12 => rom_bram_13_INIT_12,
    INIT_13 => rom_bram_13_INIT_13,
    INIT_14 => rom_bram_13_INIT_14,
    INIT_15 => rom_bram_13_INIT_15,
    INIT_16 => rom_bram_13_INIT_16,
    INIT_17 => rom_bram_13_INIT_17,
    INIT_18 => rom_bram_13_INIT_18,
    INIT_19 => rom_bram_13_INIT_19,
    INIT_1A => rom_bram_13_INIT_1A,
    INIT_1B => rom_bram_13_INIT_1B,
    INIT_1C => rom_bram_13_INIT_1C,
    INIT_1D => rom_bram_13_INIT_1D,
    INIT_1E => rom_bram_13_INIT_1E,
    INIT_1F => rom_bram_13_INIT_1F,
    INIT_20 => rom_bram_13_INIT_20,
    INIT_21 => rom_bram_13_INIT_21,
    INIT_22 => rom_bram_13_INIT_22,
    INIT_23 => rom_bram_13_INIT_23,
    INIT_24 => rom_bram_13_INIT_24,
    INIT_25 => rom_bram_13_INIT_25,
    INIT_26 => rom_bram_13_INIT_26,
    INIT_27 => rom_bram_13_INIT_27,
    INIT_28 => rom_bram_13_INIT_28,
    INIT_29 => rom_bram_13_INIT_29,
    INIT_2A => rom_bram_13_INIT_2A,
    INIT_2B => rom_bram_13_INIT_2B,
    INIT_2C => rom_bram_13_INIT_2C,
    INIT_2D => rom_bram_13_INIT_2D,
    INIT_2E => rom_bram_13_INIT_2E,
    INIT_2F => rom_bram_13_INIT_2F,
    INIT_30 => rom_bram_13_INIT_30,
    INIT_31 => rom_bram_13_INIT_31,
    INIT_32 => rom_bram_13_INIT_32,
    INIT_33 => rom_bram_13_INIT_33,
    INIT_34 => rom_bram_13_INIT_34,
    INIT_35 => rom_bram_13_INIT_35,
    INIT_36 => rom_bram_13_INIT_36,
    INIT_37 => rom_bram_13_INIT_37,
    INIT_38 => rom_bram_13_INIT_38,
    INIT_39 => rom_bram_13_INIT_39,
    INIT_3A => rom_bram_13_INIT_3A,
    INIT_3B => rom_bram_13_INIT_3B,
    INIT_3C => rom_bram_13_INIT_3C,
    INIT_3D => rom_bram_13_INIT_3D,
    INIT_3E => rom_bram_13_INIT_3E,
    INIT_3F => rom_bram_13_INIT_3F )
  PORT MAP( 
    DO => rom_bram_13_dat_o,
    dop => OPEN,    
    di => "00000000",
    dip => "0",
    addr => adr_i(10 DOWNTO 0), 
    clk => clk_i,    
    en => '1',
    ssr => '0',
    we => '0' ); 
  
  -- BRAM 14 in address space [0x0000A000:0x0000A7FF], bit lane [7:0]
  rom_bram_14 : RAMB16_S9 
  GENERIC MAP(
    INIT_00 => rom_bram_14_INIT_00,
    INIT_01 => rom_bram_14_INIT_01,
    INIT_02 => rom_bram_14_INIT_02,
    INIT_03 => rom_bram_14_INIT_03,
    INIT_04 => rom_bram_14_INIT_04,
    INIT_05 => rom_bram_14_INIT_05,
    INIT_06 => rom_bram_14_INIT_06,
    INIT_07 => rom_bram_14_INIT_07,
    INIT_08 => rom_bram_14_INIT_08,
    INIT_09 => rom_bram_14_INIT_09,
    INIT_0A => rom_bram_14_INIT_0A,
    INIT_0B => rom_bram_14_INIT_0B,
    INIT_0C => rom_bram_14_INIT_0C,
    INIT_0D => rom_bram_14_INIT_0D,
    INIT_0E => rom_bram_14_INIT_0E,
    INIT_0F => rom_bram_14_INIT_0F,
    INIT_10 => rom_bram_14_INIT_10,
    INIT_11 => rom_bram_14_INIT_11,
    INIT_12 => rom_bram_14_INIT_12,
    INIT_13 => rom_bram_14_INIT_13,
    INIT_14 => rom_bram_14_INIT_14,
    INIT_15 => rom_bram_14_INIT_15,
    INIT_16 => rom_bram_14_INIT_16,
    INIT_17 => rom_bram_14_INIT_17,
    INIT_18 => rom_bram_14_INIT_18,
    INIT_19 => rom_bram_14_INIT_19,
    INIT_1A => rom_bram_14_INIT_1A,
    INIT_1B => rom_bram_14_INIT_1B,
    INIT_1C => rom_bram_14_INIT_1C,
    INIT_1D => rom_bram_14_INIT_1D,
    INIT_1E => rom_bram_14_INIT_1E,
    INIT_1F => rom_bram_14_INIT_1F,
    INIT_20 => rom_bram_14_INIT_20,
    INIT_21 => rom_bram_14_INIT_21,
    INIT_22 => rom_bram_14_INIT_22,
    INIT_23 => rom_bram_14_INIT_23,
    INIT_24 => rom_bram_14_INIT_24,
    INIT_25 => rom_bram_14_INIT_25,
    INIT_26 => rom_bram_14_INIT_26,
    INIT_27 => rom_bram_14_INIT_27,
    INIT_28 => rom_bram_14_INIT_28,
    INIT_29 => rom_bram_14_INIT_29,
    INIT_2A => rom_bram_14_INIT_2A,
    INIT_2B => rom_bram_14_INIT_2B,
    INIT_2C => rom_bram_14_INIT_2C,
    INIT_2D => rom_bram_14_INIT_2D,
    INIT_2E => rom_bram_14_INIT_2E,
    INIT_2F => rom_bram_14_INIT_2F,
    INIT_30 => rom_bram_14_INIT_30,
    INIT_31 => rom_bram_14_INIT_31,
    INIT_32 => rom_bram_14_INIT_32,
    INIT_33 => rom_bram_14_INIT_33,
    INIT_34 => rom_bram_14_INIT_34,
    INIT_35 => rom_bram_14_INIT_35,
    INIT_36 => rom_bram_14_INIT_36,
    INIT_37 => rom_bram_14_INIT_37,
    INIT_38 => rom_bram_14_INIT_38,
    INIT_39 => rom_bram_14_INIT_39,
    INIT_3A => rom_bram_14_INIT_3A,
    INIT_3B => rom_bram_14_INIT_3B,
    INIT_3C => rom_bram_14_INIT_3C,
    INIT_3D => rom_bram_14_INIT_3D,
    INIT_3E => rom_bram_14_INIT_3E,
    INIT_3F => rom_bram_14_INIT_3F )
  PORT MAP( 
    DO => rom_bram_14_dat_o,
    dop => OPEN,    
    di => "00000000",
    dip => "0",
    addr => adr_i(10 DOWNTO 0), 
    clk => clk_i,    
    en => '1',
    ssr => '0',
    we => '0' );

  -- BRAM 15 in address space [0x0000A800:0x0000AFFF], bit lane [7:0]
  rom_bram_15 : RAMB16_S9 
  GENERIC MAP(
    INIT_00 => rom_bram_15_INIT_00,
    INIT_01 => rom_bram_15_INIT_01,
    INIT_02 => rom_bram_15_INIT_02,
    INIT_03 => rom_bram_15_INIT_03,
    INIT_04 => rom_bram_15_INIT_04,
    INIT_05 => rom_bram_15_INIT_05,
    INIT_06 => rom_bram_15_INIT_06,
    INIT_07 => rom_bram_15_INIT_07,
    INIT_08 => rom_bram_15_INIT_08,
    INIT_09 => rom_bram_15_INIT_09,
    INIT_0A => rom_bram_15_INIT_0A,
    INIT_0B => rom_bram_15_INIT_0B,
    INIT_0C => rom_bram_15_INIT_0C,
    INIT_0D => rom_bram_15_INIT_0D,
    INIT_0E => rom_bram_15_INIT_0E,
    INIT_0F => rom_bram_15_INIT_0F,
    INIT_10 => rom_bram_15_INIT_10,
    INIT_11 => rom_bram_15_INIT_11,
    INIT_12 => rom_bram_15_INIT_12,
    INIT_13 => rom_bram_15_INIT_13,
    INIT_14 => rom_bram_15_INIT_14,
    INIT_15 => rom_bram_15_INIT_15,
    INIT_16 => rom_bram_15_INIT_16,
    INIT_17 => rom_bram_15_INIT_17,
    INIT_18 => rom_bram_15_INIT_18,
    INIT_19 => rom_bram_15_INIT_19,
    INIT_1A => rom_bram_15_INIT_1A,
    INIT_1B => rom_bram_15_INIT_1B,
    INIT_1C => rom_bram_15_INIT_1C,
    INIT_1D => rom_bram_15_INIT_1D,
    INIT_1E => rom_bram_15_INIT_1E,
    INIT_1F => rom_bram_15_INIT_1F,
    INIT_20 => rom_bram_15_INIT_20,
    INIT_21 => rom_bram_15_INIT_21,
    INIT_22 => rom_bram_15_INIT_22,
    INIT_23 => rom_bram_15_INIT_23,
    INIT_24 => rom_bram_15_INIT_24,
    INIT_25 => rom_bram_15_INIT_25,
    INIT_26 => rom_bram_15_INIT_26,
    INIT_27 => rom_bram_15_INIT_27,
    INIT_28 => rom_bram_15_INIT_28,
    INIT_29 => rom_bram_15_INIT_29,
    INIT_2A => rom_bram_15_INIT_2A,
    INIT_2B => rom_bram_15_INIT_2B,
    INIT_2C => rom_bram_15_INIT_2C,
    INIT_2D => rom_bram_15_INIT_2D,
    INIT_2E => rom_bram_15_INIT_2E,
    INIT_2F => rom_bram_15_INIT_2F,
    INIT_30 => rom_bram_15_INIT_30,
    INIT_31 => rom_bram_15_INIT_31,
    INIT_32 => rom_bram_15_INIT_32,
    INIT_33 => rom_bram_15_INIT_33,
    INIT_34 => rom_bram_15_INIT_34,
    INIT_35 => rom_bram_15_INIT_35,
    INIT_36 => rom_bram_15_INIT_36,
    INIT_37 => rom_bram_15_INIT_37,
    INIT_38 => rom_bram_15_INIT_38,
    INIT_39 => rom_bram_15_INIT_39,
    INIT_3A => rom_bram_15_INIT_3A,
    INIT_3B => rom_bram_15_INIT_3B,
    INIT_3C => rom_bram_15_INIT_3C,
    INIT_3D => rom_bram_15_INIT_3D,
    INIT_3E => rom_bram_15_INIT_3E,
    INIT_3F => rom_bram_15_INIT_3F )
  PORT MAP( 
    DO => rom_bram_15_dat_o,
    dop => OPEN,    
    di => "00000000",
    dip => "0",
    addr => adr_i(10 DOWNTO 0), 
    clk => clk_i,    
    en => '1',
    ssr => '0',
    we => '0' );
    
  -- BRAM 16 in address space [0x0000B000:0x0000B7FF], bit lane [7:0]
  rom_bram_16 : RAMB16_S9 
  GENERIC MAP(
    INIT_00 => rom_bram_16_INIT_00,
    INIT_01 => rom_bram_16_INIT_01,
    INIT_02 => rom_bram_16_INIT_02,
    INIT_03 => rom_bram_16_INIT_03,
    INIT_04 => rom_bram_16_INIT_04,
    INIT_05 => rom_bram_16_INIT_05,
    INIT_06 => rom_bram_16_INIT_06,
    INIT_07 => rom_bram_16_INIT_07,
    INIT_08 => rom_bram_16_INIT_08,
    INIT_09 => rom_bram_16_INIT_09,
    INIT_0A => rom_bram_16_INIT_0A,
    INIT_0B => rom_bram_16_INIT_0B,
    INIT_0C => rom_bram_16_INIT_0C,
    INIT_0D => rom_bram_16_INIT_0D,
    INIT_0E => rom_bram_16_INIT_0E,
    INIT_0F => rom_bram_16_INIT_0F,
    INIT_10 => rom_bram_16_INIT_10,
    INIT_11 => rom_bram_16_INIT_11,
    INIT_12 => rom_bram_16_INIT_12,
    INIT_13 => rom_bram_16_INIT_13,
    INIT_14 => rom_bram_16_INIT_14,
    INIT_15 => rom_bram_16_INIT_15,
    INIT_16 => rom_bram_16_INIT_16,
    INIT_17 => rom_bram_16_INIT_17,
    INIT_18 => rom_bram_16_INIT_18,
    INIT_19 => rom_bram_16_INIT_19,
    INIT_1A => rom_bram_16_INIT_1A,
    INIT_1B => rom_bram_16_INIT_1B,
    INIT_1C => rom_bram_16_INIT_1C,
    INIT_1D => rom_bram_16_INIT_1D,
    INIT_1E => rom_bram_16_INIT_1E,
    INIT_1F => rom_bram_16_INIT_1F,
    INIT_20 => rom_bram_16_INIT_20,
    INIT_21 => rom_bram_16_INIT_21,
    INIT_22 => rom_bram_16_INIT_22,
    INIT_23 => rom_bram_16_INIT_23,
    INIT_24 => rom_bram_16_INIT_24,
    INIT_25 => rom_bram_16_INIT_25,
    INIT_26 => rom_bram_16_INIT_26,
    INIT_27 => rom_bram_16_INIT_27,
    INIT_28 => rom_bram_16_INIT_28,
    INIT_29 => rom_bram_16_INIT_29,
    INIT_2A => rom_bram_16_INIT_2A,
    INIT_2B => rom_bram_16_INIT_2B,
    INIT_2C => rom_bram_16_INIT_2C,
    INIT_2D => rom_bram_16_INIT_2D,
    INIT_2E => rom_bram_16_INIT_2E,
    INIT_2F => rom_bram_16_INIT_2F,
    INIT_30 => rom_bram_16_INIT_30,
    INIT_31 => rom_bram_16_INIT_31,
    INIT_32 => rom_bram_16_INIT_32,
    INIT_33 => rom_bram_16_INIT_33,
    INIT_34 => rom_bram_16_INIT_34,
    INIT_35 => rom_bram_16_INIT_35,
    INIT_36 => rom_bram_16_INIT_36,
    INIT_37 => rom_bram_16_INIT_37,
    INIT_38 => rom_bram_16_INIT_38,
    INIT_39 => rom_bram_16_INIT_39,
    INIT_3A => rom_bram_16_INIT_3A,
    INIT_3B => rom_bram_16_INIT_3B,
    INIT_3C => rom_bram_16_INIT_3C,
    INIT_3D => rom_bram_16_INIT_3D,
    INIT_3E => rom_bram_16_INIT_3E,
    INIT_3F => rom_bram_16_INIT_3F )
  PORT MAP( 
    DO => rom_bram_16_dat_o,
    dop => OPEN,    
    di => "00000000",
    dip => "0",
    addr => adr_i(10 DOWNTO 0), 
    clk => clk_i,    
    en => '1',
    ssr => '0',
    we => '0' );
    
  -- BRAM 17 in address space [0x0000B800:0x0000BFFF], bit lane [7:0]
  rom_bram_17 : RAMB16_S9 
  GENERIC MAP(
    INIT_00 => rom_bram_17_INIT_00,
    INIT_01 => rom_bram_17_INIT_01,
    INIT_02 => rom_bram_17_INIT_02,
    INIT_03 => rom_bram_17_INIT_03,
    INIT_04 => rom_bram_17_INIT_04,
    INIT_05 => rom_bram_17_INIT_05,
    INIT_06 => rom_bram_17_INIT_06,
    INIT_07 => rom_bram_17_INIT_07,
    INIT_08 => rom_bram_17_INIT_08,
    INIT_09 => rom_bram_17_INIT_09,
    INIT_0A => rom_bram_17_INIT_0A,
    INIT_0B => rom_bram_17_INIT_0B,
    INIT_0C => rom_bram_17_INIT_0C,
    INIT_0D => rom_bram_17_INIT_0D,
    INIT_0E => rom_bram_17_INIT_0E,
    INIT_0F => rom_bram_17_INIT_0F,
    INIT_10 => rom_bram_17_INIT_10,
    INIT_11 => rom_bram_17_INIT_11,
    INIT_12 => rom_bram_17_INIT_12,
    INIT_13 => rom_bram_17_INIT_13,
    INIT_14 => rom_bram_17_INIT_14,
    INIT_15 => rom_bram_17_INIT_15,
    INIT_16 => rom_bram_17_INIT_16,
    INIT_17 => rom_bram_17_INIT_17,
    INIT_18 => rom_bram_17_INIT_18,
    INIT_19 => rom_bram_17_INIT_19,
    INIT_1A => rom_bram_17_INIT_1A,
    INIT_1B => rom_bram_17_INIT_1B,
    INIT_1C => rom_bram_17_INIT_1C,
    INIT_1D => rom_bram_17_INIT_1D,
    INIT_1E => rom_bram_17_INIT_1E,
    INIT_1F => rom_bram_17_INIT_1F,
    INIT_20 => rom_bram_17_INIT_20,
    INIT_21 => rom_bram_17_INIT_21,
    INIT_22 => rom_bram_17_INIT_22,
    INIT_23 => rom_bram_17_INIT_23,
    INIT_24 => rom_bram_17_INIT_24,
    INIT_25 => rom_bram_17_INIT_25,
    INIT_26 => rom_bram_17_INIT_26,
    INIT_27 => rom_bram_17_INIT_27,
    INIT_28 => rom_bram_17_INIT_28,
    INIT_29 => rom_bram_17_INIT_29,
    INIT_2A => rom_bram_17_INIT_2A,
    INIT_2B => rom_bram_17_INIT_2B,
    INIT_2C => rom_bram_17_INIT_2C,
    INIT_2D => rom_bram_17_INIT_2D,
    INIT_2E => rom_bram_17_INIT_2E,
    INIT_2F => rom_bram_17_INIT_2F,
    INIT_30 => rom_bram_17_INIT_30,
    INIT_31 => rom_bram_17_INIT_31,
    INIT_32 => rom_bram_17_INIT_32,
    INIT_33 => rom_bram_17_INIT_33,
    INIT_34 => rom_bram_17_INIT_34,
    INIT_35 => rom_bram_17_INIT_35,
    INIT_36 => rom_bram_17_INIT_36,
    INIT_37 => rom_bram_17_INIT_37,
    INIT_38 => rom_bram_17_INIT_38,
    INIT_39 => rom_bram_17_INIT_39,
    INIT_3A => rom_bram_17_INIT_3A,
    INIT_3B => rom_bram_17_INIT_3B,
    INIT_3C => rom_bram_17_INIT_3C,
    INIT_3D => rom_bram_17_INIT_3D,
    INIT_3E => rom_bram_17_INIT_3E,
    INIT_3F => rom_bram_17_INIT_3F )
  PORT MAP( 
    DO => rom_bram_17_dat_o,
    dop => OPEN,    
    di => "00000000",
    dip => "0",
    addr => adr_i(10 DOWNTO 0), 
    clk => clk_i,    
    en => '1',
    ssr => '0',
    we => '0' );

  -- BRAM 18 in address space [0x0000C000:0x0000C7FF], bit lane [7:0]
  rom_bram_18 : RAMB16_S9 
  GENERIC MAP(
    INIT_00 => rom_bram_18_INIT_00,
    INIT_01 => rom_bram_18_INIT_01,
    INIT_02 => rom_bram_18_INIT_02,
    INIT_03 => rom_bram_18_INIT_03,
    INIT_04 => rom_bram_18_INIT_04,
    INIT_05 => rom_bram_18_INIT_05,
    INIT_06 => rom_bram_18_INIT_06,
    INIT_07 => rom_bram_18_INIT_07,
    INIT_08 => rom_bram_18_INIT_08,
    INIT_09 => rom_bram_18_INIT_09,
    INIT_0A => rom_bram_18_INIT_0A,
    INIT_0B => rom_bram_18_INIT_0B,
    INIT_0C => rom_bram_18_INIT_0C,
    INIT_0D => rom_bram_18_INIT_0D,
    INIT_0E => rom_bram_18_INIT_0E,
    INIT_0F => rom_bram_18_INIT_0F,
    INIT_10 => rom_bram_18_INIT_10,
    INIT_11 => rom_bram_18_INIT_11,
    INIT_12 => rom_bram_18_INIT_12,
    INIT_13 => rom_bram_18_INIT_13,
    INIT_14 => rom_bram_18_INIT_14,
    INIT_15 => rom_bram_18_INIT_15,
    INIT_16 => rom_bram_18_INIT_16,
    INIT_17 => rom_bram_18_INIT_17,
    INIT_18 => rom_bram_18_INIT_18,
    INIT_19 => rom_bram_18_INIT_19,
    INIT_1A => rom_bram_18_INIT_1A,
    INIT_1B => rom_bram_18_INIT_1B,
    INIT_1C => rom_bram_18_INIT_1C,
    INIT_1D => rom_bram_18_INIT_1D,
    INIT_1E => rom_bram_18_INIT_1E,
    INIT_1F => rom_bram_18_INIT_1F,
    INIT_20 => rom_bram_18_INIT_20,
    INIT_21 => rom_bram_18_INIT_21,
    INIT_22 => rom_bram_18_INIT_22,
    INIT_23 => rom_bram_18_INIT_23,
    INIT_24 => rom_bram_18_INIT_24,
    INIT_25 => rom_bram_18_INIT_25,
    INIT_26 => rom_bram_18_INIT_26,
    INIT_27 => rom_bram_18_INIT_27,
    INIT_28 => rom_bram_18_INIT_28,
    INIT_29 => rom_bram_18_INIT_29,
    INIT_2A => rom_bram_18_INIT_2A,
    INIT_2B => rom_bram_18_INIT_2B,
    INIT_2C => rom_bram_18_INIT_2C,
    INIT_2D => rom_bram_18_INIT_2D,
    INIT_2E => rom_bram_18_INIT_2E,
    INIT_2F => rom_bram_18_INIT_2F,
    INIT_30 => rom_bram_18_INIT_30,
    INIT_31 => rom_bram_18_INIT_31,
    INIT_32 => rom_bram_18_INIT_32,
    INIT_33 => rom_bram_18_INIT_33,
    INIT_34 => rom_bram_18_INIT_34,
    INIT_35 => rom_bram_18_INIT_35,
    INIT_36 => rom_bram_18_INIT_36,
    INIT_37 => rom_bram_18_INIT_37,
    INIT_38 => rom_bram_18_INIT_38,
    INIT_39 => rom_bram_18_INIT_39,
    INIT_3A => rom_bram_18_INIT_3A,
    INIT_3B => rom_bram_18_INIT_3B,
    INIT_3C => rom_bram_18_INIT_3C,
    INIT_3D => rom_bram_18_INIT_3D,
    INIT_3E => rom_bram_18_INIT_3E,
    INIT_3F => rom_bram_18_INIT_3F )
  PORT MAP( 
    DO => rom_bram_18_dat_o,
    dop => OPEN,    
    di => "00000000",
    dip => "0",
    addr => adr_i(10 DOWNTO 0), 
    clk => clk_i,    
    en => '1',
    ssr => '0',
    we => '0' );

  -- BRAM 19 in address space [0x0000C800:0x0000CFFF], bit lane [7:0]
  rom_bram_19 : RAMB16_S9 
  GENERIC MAP(
    INIT_00 => rom_bram_19_INIT_00,
    INIT_01 => rom_bram_19_INIT_01,
    INIT_02 => rom_bram_19_INIT_02,
    INIT_03 => rom_bram_19_INIT_03,
    INIT_04 => rom_bram_19_INIT_04,
    INIT_05 => rom_bram_19_INIT_05,
    INIT_06 => rom_bram_19_INIT_06,
    INIT_07 => rom_bram_19_INIT_07,
    INIT_08 => rom_bram_19_INIT_08,
    INIT_09 => rom_bram_19_INIT_09,
    INIT_0A => rom_bram_19_INIT_0A,
    INIT_0B => rom_bram_19_INIT_0B,
    INIT_0C => rom_bram_19_INIT_0C,
    INIT_0D => rom_bram_19_INIT_0D,
    INIT_0E => rom_bram_19_INIT_0E,
    INIT_0F => rom_bram_19_INIT_0F,
    INIT_10 => rom_bram_19_INIT_10,
    INIT_11 => rom_bram_19_INIT_11,
    INIT_12 => rom_bram_19_INIT_12,
    INIT_13 => rom_bram_19_INIT_13,
    INIT_14 => rom_bram_19_INIT_14,
    INIT_15 => rom_bram_19_INIT_15,
    INIT_16 => rom_bram_19_INIT_16,
    INIT_17 => rom_bram_19_INIT_17,
    INIT_18 => rom_bram_19_INIT_18,
    INIT_19 => rom_bram_19_INIT_19,
    INIT_1A => rom_bram_19_INIT_1A,
    INIT_1B => rom_bram_19_INIT_1B,
    INIT_1C => rom_bram_19_INIT_1C,
    INIT_1D => rom_bram_19_INIT_1D,
    INIT_1E => rom_bram_19_INIT_1E,
    INIT_1F => rom_bram_19_INIT_1F,
    INIT_20 => rom_bram_19_INIT_20,
    INIT_21 => rom_bram_19_INIT_21,
    INIT_22 => rom_bram_19_INIT_22,
    INIT_23 => rom_bram_19_INIT_23,
    INIT_24 => rom_bram_19_INIT_24,
    INIT_25 => rom_bram_19_INIT_25,
    INIT_26 => rom_bram_19_INIT_26,
    INIT_27 => rom_bram_19_INIT_27,
    INIT_28 => rom_bram_19_INIT_28,
    INIT_29 => rom_bram_19_INIT_29,
    INIT_2A => rom_bram_19_INIT_2A,
    INIT_2B => rom_bram_19_INIT_2B,
    INIT_2C => rom_bram_19_INIT_2C,
    INIT_2D => rom_bram_19_INIT_2D,
    INIT_2E => rom_bram_19_INIT_2E,
    INIT_2F => rom_bram_19_INIT_2F,
    INIT_30 => rom_bram_19_INIT_30,
    INIT_31 => rom_bram_19_INIT_31,
    INIT_32 => rom_bram_19_INIT_32,
    INIT_33 => rom_bram_19_INIT_33,
    INIT_34 => rom_bram_19_INIT_34,
    INIT_35 => rom_bram_19_INIT_35,
    INIT_36 => rom_bram_19_INIT_36,
    INIT_37 => rom_bram_19_INIT_37,
    INIT_38 => rom_bram_19_INIT_38,
    INIT_39 => rom_bram_19_INIT_39,
    INIT_3A => rom_bram_19_INIT_3A,
    INIT_3B => rom_bram_19_INIT_3B,
    INIT_3C => rom_bram_19_INIT_3C,
    INIT_3D => rom_bram_19_INIT_3D,
    INIT_3E => rom_bram_19_INIT_3E,
    INIT_3F => rom_bram_19_INIT_3F )
  PORT MAP( 
    DO => rom_bram_19_dat_o,
    dop => OPEN,    
    di => "00000000",
    dip => "0",
    addr => adr_i(10 DOWNTO 0), 
    clk => clk_i,    
    en => '1',
    ssr => '0',
    we => '0' );
    
  -- BRAM 1A in address space [0x0000D000:0x0000D7FF], bit lane [7:0]
  rom_bram_1A : RAMB16_S9 
  GENERIC MAP(
    INIT_00 => rom_bram_1A_INIT_00,
    INIT_01 => rom_bram_1A_INIT_01,
    INIT_02 => rom_bram_1A_INIT_02,
    INIT_03 => rom_bram_1A_INIT_03,
    INIT_04 => rom_bram_1A_INIT_04,
    INIT_05 => rom_bram_1A_INIT_05,
    INIT_06 => rom_bram_1A_INIT_06,
    INIT_07 => rom_bram_1A_INIT_07,
    INIT_08 => rom_bram_1A_INIT_08,
    INIT_09 => rom_bram_1A_INIT_09,
    INIT_0A => rom_bram_1A_INIT_0A,
    INIT_0B => rom_bram_1A_INIT_0B,
    INIT_0C => rom_bram_1A_INIT_0C,
    INIT_0D => rom_bram_1A_INIT_0D,
    INIT_0E => rom_bram_1A_INIT_0E,
    INIT_0F => rom_bram_1A_INIT_0F,
    INIT_10 => rom_bram_1A_INIT_10,
    INIT_11 => rom_bram_1A_INIT_11,
    INIT_12 => rom_bram_1A_INIT_12,
    INIT_13 => rom_bram_1A_INIT_13,
    INIT_14 => rom_bram_1A_INIT_14,
    INIT_15 => rom_bram_1A_INIT_15,
    INIT_16 => rom_bram_1A_INIT_16,
    INIT_17 => rom_bram_1A_INIT_17,
    INIT_18 => rom_bram_1A_INIT_18,
    INIT_19 => rom_bram_1A_INIT_19,
    INIT_1A => rom_bram_1A_INIT_1A,
    INIT_1B => rom_bram_1A_INIT_1B,
    INIT_1C => rom_bram_1A_INIT_1C,
    INIT_1D => rom_bram_1A_INIT_1D,
    INIT_1E => rom_bram_1A_INIT_1E,
    INIT_1F => rom_bram_1A_INIT_1F,
    INIT_20 => rom_bram_1A_INIT_20,
    INIT_21 => rom_bram_1A_INIT_21,
    INIT_22 => rom_bram_1A_INIT_22,
    INIT_23 => rom_bram_1A_INIT_23,
    INIT_24 => rom_bram_1A_INIT_24,
    INIT_25 => rom_bram_1A_INIT_25,
    INIT_26 => rom_bram_1A_INIT_26,
    INIT_27 => rom_bram_1A_INIT_27,
    INIT_28 => rom_bram_1A_INIT_28,
    INIT_29 => rom_bram_1A_INIT_29,
    INIT_2A => rom_bram_1A_INIT_2A,
    INIT_2B => rom_bram_1A_INIT_2B,
    INIT_2C => rom_bram_1A_INIT_2C,
    INIT_2D => rom_bram_1A_INIT_2D,
    INIT_2E => rom_bram_1A_INIT_2E,
    INIT_2F => rom_bram_1A_INIT_2F,
    INIT_30 => rom_bram_1A_INIT_30,
    INIT_31 => rom_bram_1A_INIT_31,
    INIT_32 => rom_bram_1A_INIT_32,
    INIT_33 => rom_bram_1A_INIT_33,
    INIT_34 => rom_bram_1A_INIT_34,
    INIT_35 => rom_bram_1A_INIT_35,
    INIT_36 => rom_bram_1A_INIT_36,
    INIT_37 => rom_bram_1A_INIT_37,
    INIT_38 => rom_bram_1A_INIT_38,
    INIT_39 => rom_bram_1A_INIT_39,
    INIT_3A => rom_bram_1A_INIT_3A,
    INIT_3B => rom_bram_1A_INIT_3B,
    INIT_3C => rom_bram_1A_INIT_3C,
    INIT_3D => rom_bram_1A_INIT_3D,
    INIT_3E => rom_bram_1A_INIT_3E,
    INIT_3F => rom_bram_1A_INIT_3F )
  PORT MAP( 
    DO => rom_bram_1A_dat_o,
    dop => OPEN,    
    di => "00000000",
    dip => "0",
    addr => adr_i(10 DOWNTO 0), 
    clk => clk_i,    
    en => '1',
    ssr => '0',
    we => '0' );
    
  -- BRAM 1B in address space [0x0000D800:0x0000DFFF], bit lane [7:0]
  rom_bram_1B : RAMB16_S9 
  GENERIC MAP(
    INIT_00 => rom_bram_1B_INIT_00,
    INIT_01 => rom_bram_1B_INIT_01,
    INIT_02 => rom_bram_1B_INIT_02,
    INIT_03 => rom_bram_1B_INIT_03,
    INIT_04 => rom_bram_1B_INIT_04,
    INIT_05 => rom_bram_1B_INIT_05,
    INIT_06 => rom_bram_1B_INIT_06,
    INIT_07 => rom_bram_1B_INIT_07,
    INIT_08 => rom_bram_1B_INIT_08,
    INIT_09 => rom_bram_1B_INIT_09,
    INIT_0A => rom_bram_1B_INIT_0A,
    INIT_0B => rom_bram_1B_INIT_0B,
    INIT_0C => rom_bram_1B_INIT_0C,
    INIT_0D => rom_bram_1B_INIT_0D,
    INIT_0E => rom_bram_1B_INIT_0E,
    INIT_0F => rom_bram_1B_INIT_0F,
    INIT_10 => rom_bram_1B_INIT_10,
    INIT_11 => rom_bram_1B_INIT_11,
    INIT_12 => rom_bram_1B_INIT_12,
    INIT_13 => rom_bram_1B_INIT_13,
    INIT_14 => rom_bram_1B_INIT_14,
    INIT_15 => rom_bram_1B_INIT_15,
    INIT_16 => rom_bram_1B_INIT_16,
    INIT_17 => rom_bram_1B_INIT_17,
    INIT_18 => rom_bram_1B_INIT_18,
    INIT_19 => rom_bram_1B_INIT_19,
    INIT_1A => rom_bram_1B_INIT_1A,
    INIT_1B => rom_bram_1B_INIT_1B,
    INIT_1C => rom_bram_1B_INIT_1C,
    INIT_1D => rom_bram_1B_INIT_1D,
    INIT_1E => rom_bram_1B_INIT_1E,
    INIT_1F => rom_bram_1B_INIT_1F,
    INIT_20 => rom_bram_1B_INIT_20,
    INIT_21 => rom_bram_1B_INIT_21,
    INIT_22 => rom_bram_1B_INIT_22,
    INIT_23 => rom_bram_1B_INIT_23,
    INIT_24 => rom_bram_1B_INIT_24,
    INIT_25 => rom_bram_1B_INIT_25,
    INIT_26 => rom_bram_1B_INIT_26,
    INIT_27 => rom_bram_1B_INIT_27,
    INIT_28 => rom_bram_1B_INIT_28,
    INIT_29 => rom_bram_1B_INIT_29,
    INIT_2A => rom_bram_1B_INIT_2A,
    INIT_2B => rom_bram_1B_INIT_2B,
    INIT_2C => rom_bram_1B_INIT_2C,
    INIT_2D => rom_bram_1B_INIT_2D,
    INIT_2E => rom_bram_1B_INIT_2E,
    INIT_2F => rom_bram_1B_INIT_2F,
    INIT_30 => rom_bram_1B_INIT_30,
    INIT_31 => rom_bram_1B_INIT_31,
    INIT_32 => rom_bram_1B_INIT_32,
    INIT_33 => rom_bram_1B_INIT_33,
    INIT_34 => rom_bram_1B_INIT_34,
    INIT_35 => rom_bram_1B_INIT_35,
    INIT_36 => rom_bram_1B_INIT_36,
    INIT_37 => rom_bram_1B_INIT_37,
    INIT_38 => rom_bram_1B_INIT_38,
    INIT_39 => rom_bram_1B_INIT_39,
    INIT_3A => rom_bram_1B_INIT_3A,
    INIT_3B => rom_bram_1B_INIT_3B,
    INIT_3C => rom_bram_1B_INIT_3C,
    INIT_3D => rom_bram_1B_INIT_3D,
    INIT_3E => rom_bram_1B_INIT_3E,
    INIT_3F => rom_bram_1B_INIT_3F )
  PORT MAP( 
    DO => rom_bram_1B_dat_o,
    dop => OPEN,    
    di => "00000000",
    dip => "0",
    addr => adr_i(10 DOWNTO 0), 
    clk => clk_i,    
    en => '1',
    ssr => '0',
    we => '0' ); 
  
  -- BRAM 1C in address space [0x0000E000:0x0000E7FF], bit lane [7:0]
  rom_bram_1C : RAMB16_S9 
  GENERIC MAP(
    INIT_00 => rom_bram_1C_INIT_00,
    INIT_01 => rom_bram_1C_INIT_01,
    INIT_02 => rom_bram_1C_INIT_02,
    INIT_03 => rom_bram_1C_INIT_03,
    INIT_04 => rom_bram_1C_INIT_04,
    INIT_05 => rom_bram_1C_INIT_05,
    INIT_06 => rom_bram_1C_INIT_06,
    INIT_07 => rom_bram_1C_INIT_07,
    INIT_08 => rom_bram_1C_INIT_08,
    INIT_09 => rom_bram_1C_INIT_09,
    INIT_0A => rom_bram_1C_INIT_0A,
    INIT_0B => rom_bram_1C_INIT_0B,
    INIT_0C => rom_bram_1C_INIT_0C,
    INIT_0D => rom_bram_1C_INIT_0D,
    INIT_0E => rom_bram_1C_INIT_0E,
    INIT_0F => rom_bram_1C_INIT_0F,
    INIT_10 => rom_bram_1C_INIT_10,
    INIT_11 => rom_bram_1C_INIT_11,
    INIT_12 => rom_bram_1C_INIT_12,
    INIT_13 => rom_bram_1C_INIT_13,
    INIT_14 => rom_bram_1C_INIT_14,
    INIT_15 => rom_bram_1C_INIT_15,
    INIT_16 => rom_bram_1C_INIT_16,
    INIT_17 => rom_bram_1C_INIT_17,
    INIT_18 => rom_bram_1C_INIT_18,
    INIT_19 => rom_bram_1C_INIT_19,
    INIT_1A => rom_bram_1C_INIT_1A,
    INIT_1B => rom_bram_1C_INIT_1B,
    INIT_1C => rom_bram_1C_INIT_1C,
    INIT_1D => rom_bram_1C_INIT_1D,
    INIT_1E => rom_bram_1C_INIT_1E,
    INIT_1F => rom_bram_1C_INIT_1F,
    INIT_20 => rom_bram_1C_INIT_20,
    INIT_21 => rom_bram_1C_INIT_21,
    INIT_22 => rom_bram_1C_INIT_22,
    INIT_23 => rom_bram_1C_INIT_23,
    INIT_24 => rom_bram_1C_INIT_24,
    INIT_25 => rom_bram_1C_INIT_25,
    INIT_26 => rom_bram_1C_INIT_26,
    INIT_27 => rom_bram_1C_INIT_27,
    INIT_28 => rom_bram_1C_INIT_28,
    INIT_29 => rom_bram_1C_INIT_29,
    INIT_2A => rom_bram_1C_INIT_2A,
    INIT_2B => rom_bram_1C_INIT_2B,
    INIT_2C => rom_bram_1C_INIT_2C,
    INIT_2D => rom_bram_1C_INIT_2D,
    INIT_2E => rom_bram_1C_INIT_2E,
    INIT_2F => rom_bram_1C_INIT_2F,
    INIT_30 => rom_bram_1C_INIT_30,
    INIT_31 => rom_bram_1C_INIT_31,
    INIT_32 => rom_bram_1C_INIT_32,
    INIT_33 => rom_bram_1C_INIT_33,
    INIT_34 => rom_bram_1C_INIT_34,
    INIT_35 => rom_bram_1C_INIT_35,
    INIT_36 => rom_bram_1C_INIT_36,
    INIT_37 => rom_bram_1C_INIT_37,
    INIT_38 => rom_bram_1C_INIT_38,
    INIT_39 => rom_bram_1C_INIT_39,
    INIT_3A => rom_bram_1C_INIT_3A,
    INIT_3B => rom_bram_1C_INIT_3B,
    INIT_3C => rom_bram_1C_INIT_3C,
    INIT_3D => rom_bram_1C_INIT_3D,
    INIT_3E => rom_bram_1C_INIT_3E,
    INIT_3F => rom_bram_1C_INIT_3F )
  PORT MAP( 
    DO => rom_bram_1C_dat_o,
    dop => OPEN,    
    di => "00000000",
    dip => "0",
    addr => adr_i(10 DOWNTO 0), 
    clk => clk_i,    
    en => '1',
    ssr => '0',
    we => '0' );

  -- BRAM 1D in address space [0x0000E800:0x0000EFFF], bit lane [7:0]
  rom_bram_1D : RAMB16_S9 
  GENERIC MAP(
    INIT_00 => rom_bram_1D_INIT_00,
    INIT_01 => rom_bram_1D_INIT_01,
    INIT_02 => rom_bram_1D_INIT_02,
    INIT_03 => rom_bram_1D_INIT_03,
    INIT_04 => rom_bram_1D_INIT_04,
    INIT_05 => rom_bram_1D_INIT_05,
    INIT_06 => rom_bram_1D_INIT_06,
    INIT_07 => rom_bram_1D_INIT_07,
    INIT_08 => rom_bram_1D_INIT_08,
    INIT_09 => rom_bram_1D_INIT_09,
    INIT_0A => rom_bram_1D_INIT_0A,
    INIT_0B => rom_bram_1D_INIT_0B,
    INIT_0C => rom_bram_1D_INIT_0C,
    INIT_0D => rom_bram_1D_INIT_0D,
    INIT_0E => rom_bram_1D_INIT_0E,
    INIT_0F => rom_bram_1D_INIT_0F,
    INIT_10 => rom_bram_1D_INIT_10,
    INIT_11 => rom_bram_1D_INIT_11,
    INIT_12 => rom_bram_1D_INIT_12,
    INIT_13 => rom_bram_1D_INIT_13,
    INIT_14 => rom_bram_1D_INIT_14,
    INIT_15 => rom_bram_1D_INIT_15,
    INIT_16 => rom_bram_1D_INIT_16,
    INIT_17 => rom_bram_1D_INIT_17,
    INIT_18 => rom_bram_1D_INIT_18,
    INIT_19 => rom_bram_1D_INIT_19,
    INIT_1A => rom_bram_1D_INIT_1A,
    INIT_1B => rom_bram_1D_INIT_1B,
    INIT_1C => rom_bram_1D_INIT_1C,
    INIT_1D => rom_bram_1D_INIT_1D,
    INIT_1E => rom_bram_1D_INIT_1E,
    INIT_1F => rom_bram_1D_INIT_1F,
    INIT_20 => rom_bram_1D_INIT_20,
    INIT_21 => rom_bram_1D_INIT_21,
    INIT_22 => rom_bram_1D_INIT_22,
    INIT_23 => rom_bram_1D_INIT_23,
    INIT_24 => rom_bram_1D_INIT_24,
    INIT_25 => rom_bram_1D_INIT_25,
    INIT_26 => rom_bram_1D_INIT_26,
    INIT_27 => rom_bram_1D_INIT_27,
    INIT_28 => rom_bram_1D_INIT_28,
    INIT_29 => rom_bram_1D_INIT_29,
    INIT_2A => rom_bram_1D_INIT_2A,
    INIT_2B => rom_bram_1D_INIT_2B,
    INIT_2C => rom_bram_1D_INIT_2C,
    INIT_2D => rom_bram_1D_INIT_2D,
    INIT_2E => rom_bram_1D_INIT_2E,
    INIT_2F => rom_bram_1D_INIT_2F,
    INIT_30 => rom_bram_1D_INIT_30,
    INIT_31 => rom_bram_1D_INIT_31,
    INIT_32 => rom_bram_1D_INIT_32,
    INIT_33 => rom_bram_1D_INIT_33,
    INIT_34 => rom_bram_1D_INIT_34,
    INIT_35 => rom_bram_1D_INIT_35,
    INIT_36 => rom_bram_1D_INIT_36,
    INIT_37 => rom_bram_1D_INIT_37,
    INIT_38 => rom_bram_1D_INIT_38,
    INIT_39 => rom_bram_1D_INIT_39,
    INIT_3A => rom_bram_1D_INIT_3A,
    INIT_3B => rom_bram_1D_INIT_3B,
    INIT_3C => rom_bram_1D_INIT_3C,
    INIT_3D => rom_bram_1D_INIT_3D,
    INIT_3E => rom_bram_1D_INIT_3E,
    INIT_3F => rom_bram_1D_INIT_3F )
  PORT MAP( 
    DO => rom_bram_1D_dat_o,
    dop => OPEN,    
    di => "00000000",
    dip => "0",
    addr => adr_i(10 DOWNTO 0), 
    clk => clk_i,    
    en => '1',
    ssr => '0',
    we => '0' );
    
  -- BRAM 1E in address space [0x0000F000:0x0000F7FF], bit lane [7:0]
  rom_bram_1E : RAMB16_S9 
  GENERIC MAP(
    INIT_00 => rom_bram_1E_INIT_00,
    INIT_01 => rom_bram_1E_INIT_01,
    INIT_02 => rom_bram_1E_INIT_02,
    INIT_03 => rom_bram_1E_INIT_03,
    INIT_04 => rom_bram_1E_INIT_04,
    INIT_05 => rom_bram_1E_INIT_05,
    INIT_06 => rom_bram_1E_INIT_06,
    INIT_07 => rom_bram_1E_INIT_07,
    INIT_08 => rom_bram_1E_INIT_08,
    INIT_09 => rom_bram_1E_INIT_09,
    INIT_0A => rom_bram_1E_INIT_0A,
    INIT_0B => rom_bram_1E_INIT_0B,
    INIT_0C => rom_bram_1E_INIT_0C,
    INIT_0D => rom_bram_1E_INIT_0D,
    INIT_0E => rom_bram_1E_INIT_0E,
    INIT_0F => rom_bram_1E_INIT_0F,
    INIT_10 => rom_bram_1E_INIT_10,
    INIT_11 => rom_bram_1E_INIT_11,
    INIT_12 => rom_bram_1E_INIT_12,
    INIT_13 => rom_bram_1E_INIT_13,
    INIT_14 => rom_bram_1E_INIT_14,
    INIT_15 => rom_bram_1E_INIT_15,
    INIT_16 => rom_bram_1E_INIT_16,
    INIT_17 => rom_bram_1E_INIT_17,
    INIT_18 => rom_bram_1E_INIT_18,
    INIT_19 => rom_bram_1E_INIT_19,
    INIT_1A => rom_bram_1E_INIT_1A,
    INIT_1B => rom_bram_1E_INIT_1B,
    INIT_1C => rom_bram_1E_INIT_1C,
    INIT_1D => rom_bram_1E_INIT_1D,
    INIT_1E => rom_bram_1E_INIT_1E,
    INIT_1F => rom_bram_1E_INIT_1F,
    INIT_20 => rom_bram_1E_INIT_20,
    INIT_21 => rom_bram_1E_INIT_21,
    INIT_22 => rom_bram_1E_INIT_22,
    INIT_23 => rom_bram_1E_INIT_23,
    INIT_24 => rom_bram_1E_INIT_24,
    INIT_25 => rom_bram_1E_INIT_25,
    INIT_26 => rom_bram_1E_INIT_26,
    INIT_27 => rom_bram_1E_INIT_27,
    INIT_28 => rom_bram_1E_INIT_28,
    INIT_29 => rom_bram_1E_INIT_29,
    INIT_2A => rom_bram_1E_INIT_2A,
    INIT_2B => rom_bram_1E_INIT_2B,
    INIT_2C => rom_bram_1E_INIT_2C,
    INIT_2D => rom_bram_1E_INIT_2D,
    INIT_2E => rom_bram_1E_INIT_2E,
    INIT_2F => rom_bram_1E_INIT_2F,
    INIT_30 => rom_bram_1E_INIT_30,
    INIT_31 => rom_bram_1E_INIT_31,
    INIT_32 => rom_bram_1E_INIT_32,
    INIT_33 => rom_bram_1E_INIT_33,
    INIT_34 => rom_bram_1E_INIT_34,
    INIT_35 => rom_bram_1E_INIT_35,
    INIT_36 => rom_bram_1E_INIT_36,
    INIT_37 => rom_bram_1E_INIT_37,
    INIT_38 => rom_bram_1E_INIT_38,
    INIT_39 => rom_bram_1E_INIT_39,
    INIT_3A => rom_bram_1E_INIT_3A,
    INIT_3B => rom_bram_1E_INIT_3B,
    INIT_3C => rom_bram_1E_INIT_3C,
    INIT_3D => rom_bram_1E_INIT_3D,
    INIT_3E => rom_bram_1E_INIT_3E,
    INIT_3F => rom_bram_1E_INIT_3F )
  PORT MAP( 
    DO => rom_bram_1E_dat_o,
    dop => OPEN,    
    di => "00000000",
    dip => "0",
    addr => adr_i(10 DOWNTO 0), 
    clk => clk_i,    
    en => '1',
    ssr => '0',
    we => '0' );
    
  -- BRAM 1F in address space [0x0000F800:0x0000FFFF], bit lane [7:0]
  rom_bram_1F : RAMB16_S9 
  GENERIC MAP(
    INIT_00 => rom_bram_1F_INIT_00,
    INIT_01 => rom_bram_1F_INIT_01,
    INIT_02 => rom_bram_1F_INIT_02,
    INIT_03 => rom_bram_1F_INIT_03,
    INIT_04 => rom_bram_1F_INIT_04,
    INIT_05 => rom_bram_1F_INIT_05,
    INIT_06 => rom_bram_1F_INIT_06,
    INIT_07 => rom_bram_1F_INIT_07,
    INIT_08 => rom_bram_1F_INIT_08,
    INIT_09 => rom_bram_1F_INIT_09,
    INIT_0A => rom_bram_1F_INIT_0A,
    INIT_0B => rom_bram_1F_INIT_0B,
    INIT_0C => rom_bram_1F_INIT_0C,
    INIT_0D => rom_bram_1F_INIT_0D,
    INIT_0E => rom_bram_1F_INIT_0E,
    INIT_0F => rom_bram_1F_INIT_0F,
    INIT_10 => rom_bram_1F_INIT_10,
    INIT_11 => rom_bram_1F_INIT_11,
    INIT_12 => rom_bram_1F_INIT_12,
    INIT_13 => rom_bram_1F_INIT_13,
    INIT_14 => rom_bram_1F_INIT_14,
    INIT_15 => rom_bram_1F_INIT_15,
    INIT_16 => rom_bram_1F_INIT_16,
    INIT_17 => rom_bram_1F_INIT_17,
    INIT_18 => rom_bram_1F_INIT_18,
    INIT_19 => rom_bram_1F_INIT_19,
    INIT_1A => rom_bram_1F_INIT_1A,
    INIT_1B => rom_bram_1F_INIT_1B,
    INIT_1C => rom_bram_1F_INIT_1C,
    INIT_1D => rom_bram_1F_INIT_1D,
    INIT_1E => rom_bram_1F_INIT_1E,
    INIT_1F => rom_bram_1F_INIT_1F,
    INIT_20 => rom_bram_1F_INIT_20,
    INIT_21 => rom_bram_1F_INIT_21,
    INIT_22 => rom_bram_1F_INIT_22,
    INIT_23 => rom_bram_1F_INIT_23,
    INIT_24 => rom_bram_1F_INIT_24,
    INIT_25 => rom_bram_1F_INIT_25,
    INIT_26 => rom_bram_1F_INIT_26,
    INIT_27 => rom_bram_1F_INIT_27,
    INIT_28 => rom_bram_1F_INIT_28,
    INIT_29 => rom_bram_1F_INIT_29,
    INIT_2A => rom_bram_1F_INIT_2A,
    INIT_2B => rom_bram_1F_INIT_2B,
    INIT_2C => rom_bram_1F_INIT_2C,
    INIT_2D => rom_bram_1F_INIT_2D,
    INIT_2E => rom_bram_1F_INIT_2E,
    INIT_2F => rom_bram_1F_INIT_2F,
    INIT_30 => rom_bram_1F_INIT_30,
    INIT_31 => rom_bram_1F_INIT_31,
    INIT_32 => rom_bram_1F_INIT_32,
    INIT_33 => rom_bram_1F_INIT_33,
    INIT_34 => rom_bram_1F_INIT_34,
    INIT_35 => rom_bram_1F_INIT_35,
    INIT_36 => rom_bram_1F_INIT_36,
    INIT_37 => rom_bram_1F_INIT_37,
    INIT_38 => rom_bram_1F_INIT_38,
    INIT_39 => rom_bram_1F_INIT_39,
    INIT_3A => rom_bram_1F_INIT_3A,
    INIT_3B => rom_bram_1F_INIT_3B,
    INIT_3C => rom_bram_1F_INIT_3C,
    INIT_3D => rom_bram_1F_INIT_3D,
    INIT_3E => rom_bram_1F_INIT_3E,
    INIT_3F => rom_bram_1F_INIT_3F )
  PORT MAP( 
    DO => rom_bram_1F_dat_o,
    dop => OPEN,    
    di => "00000000",
    dip => "0",
    addr => adr_i(10 DOWNTO 0), 
    clk => clk_i,    
    en => '1',
    ssr => '0',
    we => '0' );
    
END internal_rom_64K_arch;

